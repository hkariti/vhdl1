library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;

entity background is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end background;

architecture behav of background is 

constant object_X_size : integer := 640;
constant object_Y_size : integer := 480;

type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  
constant object_color: ram_array := (
(x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bb",x"bf",x"bf",x"bf",x"bf",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9f",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bb",x"bf",x"bb",x"bf",x"bf",x"bb",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bb",x"bf",x"bb",x"bf",x"df",x"bb",x"bf",x"bf",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bb",x"bb",x"9b",x"bb",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9f",x"bf",x"bf",x"bf",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"df",x"df",x"df",x"df",x"bf",x"bb",x"9b",x"bf",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"bf",x"bf",x"bb",x"9b",x"9b",x"bb",x"bf",x"df",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"df",x"df",x"df",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"df",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bb",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bf",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"df",x"df",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"bf",x"df",x"df",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bf",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"ff",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bf",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"9b",x"bf",x"df",x"bf",x"df",x"bf",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"df",x"df",x"df",x"ff",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"9b",x"bb",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"bb",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bf",x"bf",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bf",x"bf",x"df",x"df",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"9b",x"bf",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"df",x"df",x"df",x"df",x"df",x"bb",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"df",x"df",x"df",x"df",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"df",x"df",x"df",x"df",x"df",x"bf",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"9b",x"bf",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bf",x"df",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"df",x"df",x"df",x"bb",x"bf",x"9b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"bb",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9f",x"bf",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"df",x"df",x"bb",x"9b",x"7b",x"9b",x"9b",x"bb",x"df",x"df",x"df",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bb",x"bb",x"bf",x"bb",x"bb",x"bf",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bf",x"bf",x"bf",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"df",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"df",x"df",x"df",x"bf",x"bf",x"df",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"bb",x"9b",x"9b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"df",x"df",x"bf",x"bf",x"9b",x"9b",x"bb",x"bb",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"df",x"df",x"df",x"bf",x"bf",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"9b",x"9b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"bf",x"bf",x"bf",x"df",x"df",x"bf",x"df",x"df",x"bf",x"df",x"df",x"df",x"bf",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"bb",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bb",x"bf",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"9b",x"7b",x"7b",x"7b",x"bb",x"df",x"df",x"df",x"df",x"bf",x"df",x"df",x"df",x"df",x"df",x"bb",x"9b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"bb",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"9b",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"df",x"df",x"df",x"df",x"df",x"bf",x"bb",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"9b",x"9b",x"7b",x"7b",x"9b",x"bb",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bf",x"bf",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"9b",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"bb",x"bf",x"bf",x"bf",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"df",x"df",x"df",x"df",x"df",x"bf",x"bb",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"9b",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"bb",x"9b",x"bf",x"df",x"df",x"bb",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bf",x"bf",x"bb",x"bf",x"df",x"df",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"df",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"9b",x"9b",x"7b",x"7b",x"9b",x"9b",x"df",x"df",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bb",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"bb",x"df",x"df",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"9b",x"bf",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"df",x"bf",x"9b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"df",x"df",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bf",x"bf",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bf",x"bf",x"df",x"bf",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"ff",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bf",x"df",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"9b",x"bf",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"bf",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bb",x"bb",x"bb",x"bb",x"bf",x"df",x"df",x"df",x"bf",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"bf",x"bf",x"df",x"df",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"9b",x"9b",x"bb",x"bf",x"9b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9f",x"bf",x"df",x"df",x"df",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"bb",x"df",x"df",x"df",x"bb",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"bf",x"df",x"df",x"bf",x"9b",x"7b",x"9b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"bf",x"bf",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"bf",x"bb",x"bb",x"bb",x"bf",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"bf",x"bf",x"bf",x"df",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"9b",x"7b",x"7b",x"9b",x"bb",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bf",x"df",x"df",x"df",x"df",x"df",x"bb",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"ff",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"bf",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bb",x"bf",x"bf",x"bf",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"bf",x"df",x"df",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"bf",x"df",x"df",x"bf",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"ff",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"bb",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"bf",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"bb",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bf",x"bf",x"bf",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"df",x"df",x"df",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9f",x"bb",x"bf",x"9b",x"7b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"bb",x"df",x"df",x"df",x"df",x"df",x"df",x"ff",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"df",x"df",x"df",x"9b",x"7b",x"7b",x"9b",x"bf",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"df",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"9b",x"9b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"df",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"bf",x"bb",x"bb",x"bb",x"bf",x"bf",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bb",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"ff",x"ff",x"ff",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"df",x"df",x"df",x"bb",x"7b",x"9b",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"df",x"df",x"bf",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bb",x"bb",x"bf",x"bb",x"bf",x"bf",x"bb",x"bf",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bf",x"df",x"df",x"df",x"9b",x"9b",x"bb",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bb",x"bf",x"df",x"df",x"df",x"bf",x"bb",x"bf",x"df",x"df",x"df",x"df",x"df",x"bf",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"ff",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"df",x"df",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"df",x"ff",x"ff",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bf",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"7b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bf",x"ff",x"df",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"9b",x"bb",x"bb",x"bf",x"bb",x"9b",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"bb",x"bf",x"bb",x"bb",x"bf",x"bf",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"9b",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"9b",x"bb",x"9b",x"9b",x"9b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"df",x"df",x"df",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"df",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"57",x"57",x"5b",x"7b",x"9b",x"9b",x"7b",x"77",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"57",x"36",x"32",x"37",x"7b",x"7b",x"9b",x"9b",x"7b",x"77",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"0e",x"0e",x"12",x"57",x"7b",x"9b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"57",x"57",x"57",x"57",x"7b",x"7b",x"7b",x"9b",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"0e",x"0e",x"17",x"7b",x"9b",x"9b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"57",x"37",x"37",x"37",x"17",x"33",x"37",x"37",x"37",x"7b",x"9b",x"bf",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"12",x"0e",x"0e",x"0e",x"17",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"37",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"7b",x"bb",x"bb",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"12",x"0e",x"0e",x"0e",x"12",x"17",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"32",x"12",x"12",x"13",x"13",x"13",x"17",x"13",x"13",x"17",x"7b",x"bb",x"bb",x"bb",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"12",x"0e",x"0e",x"0e",x"12",x"37",x"57",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"13",x"12",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"37",x"5b",x"9b",x"bf",x"bf",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"36",x"57",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"32",x"0e",x"0e",x"12",x"12",x"37",x"37",x"7b",x"9b",x"9b",x"9b",x"9b",x"5b",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"17",x"13",x"13",x"13",x"12",x"12",x"12",x"17",x"17",x"37",x"5b",x"9b",x"bf",x"bf",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"33",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"32",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"32",x"0e",x"0e",x"12",x"32",x"37",x"37",x"37",x"5b",x"7b",x"7b",x"57",x"37",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"37",x"12",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"37",x"5b",x"5b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"32",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"57",x"12",x"0e",x"0e",x"12",x"37",x"37",x"17",x"37",x"57",x"57",x"37",x"37",x"37",x"5b",x"7b",x"5b",x"5b",x"5b",x"57",x"33",x"12",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"32",x"0e",x"0e",x"12",x"37",x"37",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"5b",x"3b",x"3b",x"37",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"df",x"ff",x"df",x"df",x"bf",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"37",x"12",x"0e",x"12",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"3b",x"17",x"12",x"17",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"0e",x"13",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"37",x"13",x"13",x"57",x"37",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"33",x"0e",x"12",x"37",x"37",x"37",x"37",x"37",x"17",x"37",x"5b",x"37",x"3b",x"3b",x"17",x"12",x"57",x"7b",x"57",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"32",x"0e",x"13",x"37",x"3b",x"37",x"37",x"37",x"5b",x"7b",x"3b",x"3b",x"37",x"13",x"37",x"7b",x"7b",x"7b",x"37",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"df",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"12",x"12",x"17",x"37",x"37",x"5b",x"5b",x"7b",x"7b",x"5b",x"37",x"13",x"13",x"5b",x"7b",x"5b",x"7b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"57",x"3b",x"37",x"57",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"33",x"57",x"7b",x"7b",x"7b",x"7b",x"7b",x"32",x"12",x"17",x"7b",x"7b",x"5b",x"7b",x"77",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"7b",x"9b",x"9f",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"0e",x"13",x"57",x"7b",x"7b",x"7b",x"7b",x"7b",x"57",x"12",x"17",x"7b",x"7b",x"7b",x"7b",x"7b",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"57",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"33",x"33",x"57",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"37",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"37",x"17",x"17",x"17",x"37",x"57",x"7b",x"7b",x"57",x"17",x"17",x"17",x"37",x"57",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"57",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"7b",x"7b",x"5b",x"7b",x"7b",x"57",x"57",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"57",x"17",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"57",x"17",x"17",x"37",x"9b",x"bf",x"bf",x"7b",x"5b",x"5b",x"17",x"17",x"17",x"17",x"37",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"df",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"32",x"12",x"32",x"33",x"37",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"37",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"17",x"17",x"7b",x"bf",x"df",x"bf",x"9b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"5b",x"7b",x"9b",x"bf",x"df",x"df",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"5b",x"7b",x"5b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"57",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"17",x"37",x"9b",x"df",x"bf",x"df",x"9b",x"5b",x"5b",x"7b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"7b",x"9b",x"bf",x"df",x"df",x"bf",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"37",x"37",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"32",x"5b",x"5b",x"57",x"36",x"12",x"12",x"13",x"13",x"33",x"57",x"57",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"37",x"37",x"bb",x"df",x"bf",x"bf",x"9b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"57",x"7b",x"7b",x"bb",x"df",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"33",x"0e",x"12",x"32",x"32",x"37",x"57",x"5b",x"57",x"0e",x"0e",x"0e",x"12",x"12",x"37",x"37",x"57",x"57",x"37",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"33",x"37",x"57",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"57",x"9b",x"bf",x"df",x"bf",x"9b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"5b",x"7b",x"7b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"0e",x"12",x"57",x"5b",x"5b",x"5b",x"5b",x"57",x"12",x"0e",x"0e",x"12",x"36",x"5b",x"7b",x"7b",x"37",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"57",x"7b",x"5b",x"7b",x"5b",x"7b",x"bf",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"bb",x"bf",x"bf",x"7b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"0e",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"0e",x"0e",x"12",x"37",x"5b",x"5b",x"5b",x"7b",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"12",x"13",x"13",x"37",x"57",x"7b",x"7b",x"5b",x"5b",x"9b",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"5b",x"57",x"57",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"57",x"5b",x"5b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"57",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"32",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"32",x"0e",x"32",x"57",x"5b",x"5b",x"5b",x"7b",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"13",x"13",x"13",x"37",x"5b",x"5b",x"7b",x"5b",x"5b",x"9b",x"bf",x"bb",x"9b",x"7b",x"5b",x"37",x"37",x"37",x"37",x"37",x"37",x"57",x"57",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"0e",x"37",x"5b",x"5b",x"5b",x"5b",x"7b",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"13",x"13",x"12",x"37",x"7b",x"5b",x"7b",x"5b",x"5b",x"7b",x"9b",x"9b",x"7b",x"5b",x"37",x"13",x"13",x"17",x"17",x"17",x"13",x"17",x"37",x"57",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bf",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"12",x"37",x"5b",x"5b",x"5b",x"5b",x"7b",x"33",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"13",x"12",x"13",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"37",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"57",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"12",x"12",x"13",x"12",x"13",x"5b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"37",x"57",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bf",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"57",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"37",x"37",x"13",x"13",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"57",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bf",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"57",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"17",x"17",x"13",x"17",x"13",x"13",x"17",x"37",x"37",x"37",x"3b",x"37",x"5b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"37",x"37",x"57",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"32",x"16",x"13",x"12",x"12",x"12",x"12",x"12",x"13",x"57",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"13",x"13",x"13",x"13",x"13",x"37",x"5b",x"7b",x"5b",x"5b",x"5b",x"3b",x"5b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"57",x"17",x"17",x"13",x"17",x"17",x"17",x"13",x"17",x"17",x"13",x"13",x"13",x"13",x"12",x"12",x"17",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"13",x"33",x"77",x"5b",x"37",x"13",x"13",x"12",x"12",x"12",x"12",x"37",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"37",x"13",x"13",x"13",x"17",x"5b",x"9b",x"9b",x"9b",x"7b",x"5b",x"3b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"37",x"13",x"13",x"13",x"17",x"13",x"13",x"37",x"57",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"77",x"9b",x"9b",x"3b",x"37",x"13",x"12",x"12",x"12",x"13",x"13",x"37",x"37",x"37",x"37",x"57",x"5b",x"7b",x"57",x"13",x"13",x"17",x"57",x"9b",x"bb",x"bb",x"9b",x"9b",x"7b",x"5b",x"3b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"13",x"13",x"37",x"37",x"37",x"57",x"5b",x"7b",x"12",x"13",x"13",x"13",x"12",x"37",x"37",x"57",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"bf",x"9b",x"3b",x"3b",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"13",x"13",x"37",x"37",x"5b",x"5b",x"13",x"13",x"17",x"5b",x"bb",x"bb",x"9b",x"9b",x"bf",x"9b",x"5b",x"3b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"13",x"57",x"5b",x"7b",x"7b",x"7b",x"7b",x"12",x"13",x"13",x"13",x"37",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"9b",x"bb",x"9b",x"37",x"3b",x"12",x"12",x"12",x"37",x"13",x"13",x"13",x"12",x"13",x"13",x"12",x"12",x"37",x"7b",x"37",x"13",x"17",x"7b",x"bb",x"9b",x"9b",x"9b",x"bf",x"9b",x"5b",x"3b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"12",x"57",x"7b",x"5b",x"5b",x"5b",x"5b",x"37",x"13",x"12",x"37",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"3b",x"37",x"3b",x"37",x"37",x"57",x"57",x"37",x"12",x"12",x"13",x"13",x"13",x"37",x"37",x"5b",x"5b",x"57",x"37",x"17",x"7b",x"bb",x"9b",x"9b",x"9b",x"bb",x"9b",x"5b",x"3b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"37",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"57",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bf",x"bf",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"37",x"17",x"37",x"5b",x"5b",x"5b",x"7b",x"7b",x"57",x"12",x"12",x"13",x"13",x"37",x"57",x"5b",x"5b",x"5b",x"7b",x"37",x"37",x"5b",x"bb",x"bb",x"9b",x"9b",x"bb",x"9b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"12",x"37",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"37",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"57",x"12",x"13",x"12",x"57",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"9b",x"bb",x"9b",x"bb",x"bb",x"7b",x"3b",x"1b",x"3b",x"37",x"3b",x"37",x"12",x"12",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"32",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"12",x"12",x"37",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"3b",x"37",x"37",x"3b",x"17",x"12",x"12",x"33",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"5b",x"7b",x"9b",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"12",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"37",x"3b",x"7b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"37",x"12",x"12",x"37",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"5b",x"7b",x"bb",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"57",x"17",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"3b",x"17",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"37",x"37",x"37",x"37",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"bb",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"57",x"17",x"57",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"5b",x"3b",x"37",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"17",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"9b",x"bb",x"9b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"57",x"37",x"37",x"17",x"37",x"37",x"37",x"57",x"57",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"37",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"37",x"37",x"17",x"37",x"17",x"37",x"37",x"37",x"37",x"37",x"57",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"37",x"37",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"37",x"17",x"37",x"17",x"37",x"37",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"37",x"57",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bb",x"bb",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"df",x"df",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"12",x"12",x"12",x"12",x"33",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"ff",x"ff",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b"),
(x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"37",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"33",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"7b",x"5b",x"9b",x"df",x"ff",x"ff",x"ff",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"37",x"17",x"17",x"37",x"37",x"17",x"17",x"37",x"17",x"17",x"37",x"17",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"57",x"57",x"57",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"9b",x"df",x"ff",x"ff",x"df",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"37",x"37",x"17",x"17",x"17",x"37",x"37",x"57",x"57",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"9b",x"bf",x"ff",x"ff",x"bf",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"17",x"16",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"16",x"37",x"57",x"5b",x"5b",x"37",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"9b",x"bb",x"bb",x"9b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"16",x"17",x"17",x"17",x"17",x"5b",x"5b",x"5b",x"5b",x"57",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"13",x"37",x"57",x"5b",x"5b",x"37",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"13",x"17",x"17",x"37",x"5b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"36",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"16",x"17",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"57",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"17",x"17",x"17",x"17",x"17",x"57",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"7b",x"7b",x"57",x"37",x"17",x"17",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"37",x"37",x"17",x"16",x"17",x"17",x"17",x"17",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"12",x"12",x"12",x"12",x"12",x"13",x"16",x"13",x"17",x"17",x"17",x"17",x"37",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"7b",x"9b",x"9b",x"7b",x"3b",x"17",x"37",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"37",x"57",x"37",x"5b",x"9b",x"bb",x"9b",x"3b",x"3b",x"17",x"16",x"17",x"37",x"17",x"37",x"37",x"37",x"5b",x"7b",x"5b",x"5b",x"5b",x"33",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"37",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"9b",x"9b",x"7b",x"17",x"37",x"37",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"36",x"7b",x"bf",x"9b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"57",x"7b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"37",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"9b",x"9b",x"9b",x"9b",x"7b",x"17",x"37",x"37",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"0e",x"0e",x"32",x"57",x"7b",x"7b",x"37",x"3b",x"37",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"17",x"12",x"13",x"13",x"12",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"5b",x"9b",x"9b",x"9b",x"9b",x"9b",x"37",x"37",x"37",x"12",x"12",x"12",x"12",x"37",x"12",x"0e",x"0e",x"0e",x"12",x"37",x"57",x"37",x"37",x"3b",x"37",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"37",x"5b",x"5b",x"5b",x"7b",x"5b",x"37",x"13",x"13",x"13",x"12",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"bb",x"bb",x"bb",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"7b",x"9b",x"9b",x"9b",x"7b",x"37",x"17",x"37",x"37",x"37",x"37",x"5b",x"3b",x"12",x"0e",x"0e",x"0e",x"12",x"37",x"37",x"37",x"37",x"37",x"37",x"16",x"17",x"17",x"17",x"37",x"37",x"17",x"37",x"5b",x"7b",x"5b",x"7b",x"5b",x"57",x"13",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"bf",x"bb",x"9b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"7b",x"7b",x"9b",x"7b",x"5b",x"37",x"17",x"37",x"57",x"57",x"5b",x"5b",x"5b",x"12",x"0e",x"0e",x"0e",x"13",x"37",x"57",x"37",x"37",x"13",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"37",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"37",x"12",x"13",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"df",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"33"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"57",x"5b",x"3b",x"57",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"37",x"57",x"5b",x"5b",x"3b",x"3b",x"5b",x"37",x"0e",x"0e",x"12",x"37",x"5b",x"5b",x"37",x"12",x"12",x"12",x"37",x"17",x"17",x"17",x"37",x"37",x"17",x"37",x"57",x"5b",x"5b",x"5b",x"7b",x"7b",x"57",x"17",x"12",x"13",x"13",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"bf",x"bf",x"bf",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"57",x"37",x"12",x"0e"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"0e",x"0e",x"37",x"3b",x"3b",x"5b",x"3b",x"32",x"0e",x"12",x"13",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"57",x"5b",x"37",x"12",x"17",x"37",x"37",x"57",x"5b",x"7b",x"57",x"17",x"17",x"17",x"12",x"17",x"37",x"37",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"bb",x"bf",x"bb",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"37",x"32",x"0e",x"0e",x"0e",x"0e"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"0e",x"37",x"5b",x"3b",x"3b",x"3b",x"37",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"17",x"37",x"17",x"17",x"17",x"37",x"5b",x"57",x"37",x"12",x"57",x"5b",x"5b",x"5b",x"7b",x"57",x"17",x"17",x"13",x"17",x"37",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"37",x"32",x"12",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"32",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"0e",x"12",x"17",x"17",x"37",x"37",x"5b",x"57",x"37",x"17",x"37",x"37",x"37",x"17",x"17",x"57",x"5b",x"37",x"17",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"13",x"12",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"bb",x"bb",x"bb",x"9b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"37",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"57",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"37",x"12",x"12",x"37",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"17",x"37",x"17",x"37",x"57",x"5b",x"7b",x"7b",x"5b",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"bb",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"3b",x"5b",x"37",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"12",x"12",x"37",x"5b",x"7b",x"5b",x"5b",x"5b",x"37",x"17",x"37",x"37",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"57",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"17",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"bb",x"bb",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"37",x"3b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"37",x"32",x"37",x"5b",x"7b",x"5b",x"5b",x"7b",x"37",x"17",x"37",x"57",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"9f",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"32",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"5b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"7b",x"37",x"17",x"37",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"37",x"37",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"37",x"5b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"5b",x"5b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"1b",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"5b",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"17",x"1b",x"3b",x"3b",x"3b",x"37",x"1b",x"1b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"37",x"37",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"12",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"3b",x"5b",x"5b",x"7b",x"9b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"37",x"3b",x"1b",x"37",x"3b",x"3b",x"37",x"3b",x"37",x"17",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"1b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"9b",x"bb",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"3b",x"3b",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"37",x"37",x"37",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"37",x"17",x"1b",x"1b",x"37",x"1b",x"1b",x"1b",x"12",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"37",x"3b",x"3b",x"1b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"bb",x"bb",x"bb",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"7b",x"9b",x"bf",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"57",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"1b",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"12",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"9b",x"bb",x"9b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"bf",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"17",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"12",x"12",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"7b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"9b",x"df",x"df",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"12",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"0e",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"57",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"7b",x"9b",x"9b",x"7b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"df",x"df",x"df",x"bf",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"12",x"12",x"37",x"3b",x"37",x"3b",x"3b",x"37",x"1b",x"1b",x"3b",x"1b",x"12",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"3b",x"17",x"3b",x"1b",x"1b",x"17",x"12",x"0a",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"9b",x"df",x"df",x"df",x"bb",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"16",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"1b",x"37",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"12",x"0e",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"1b",x"1b",x"1b",x"1b",x"3b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"bb",x"df",x"df",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"12",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"37",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"3b",x"3b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"3b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"37",x"3b",x"37",x"12",x"12",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"1b",x"3b",x"37",x"12",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"37",x"37",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"1b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"12",x"12",x"12",x"0e",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"32",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"12",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"37",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"57",x"5b",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"37",x"3b",x"17",x"17",x"3b",x"1b",x"37",x"3b",x"3b",x"37",x"37",x"1b",x"37",x"3b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"0e",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"37",x"37",x"17",x"17",x"17",x"37",x"37",x"3b",x"3b",x"3b",x"17",x"37",x"3b",x"1b",x"1b",x"3b",x"3b",x"1b",x"37",x"3b",x"3b",x"37",x"12",x"0e",x"12",x"17",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"37",x"5b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"1b",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"1b",x"17",x"3b",x"3b",x"37",x"37",x"3b",x"37",x"37",x"1b",x"37",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"0e",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"37",x"37",x"37",x"37",x"3b",x"37",x"17",x"1b",x"37",x"1b",x"1b",x"37",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"37",x"3b",x"37",x"17",x"0e",x"0e",x"17",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"9b",x"9b",x"9b",x"7b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"37",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"37",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"1b",x"3b",x"37",x"32",x"12",x"17",x"1b",x"37",x"37",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"3b",x"9b",x"bb",x"9b",x"7b",x"5b",x"3b",x"17",x"3b",x"3b",x"3b",x"5b",x"9b",x"9b",x"7b",x"5b",x"7b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"1b",x"1b",x"1b",x"3b",x"37",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"37",x"37",x"3b",x"17",x"1b",x"1b",x"37",x"37",x"37",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"37",x"33",x"13",x"1b",x"1b",x"17",x"37",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"3b",x"7b",x"9b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"7b",x"bb",x"bb",x"9b",x"7b",x"7b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"37",x"17",x"3b",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"3b",x"3b",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"0e",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"1b",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"37",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"13",x"3b",x"1b",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"3b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"7b",x"9b",x"bb",x"bb",x"9b",x"9b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"3b",x"17",x"12",x"13",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"0e",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"13",x"1b",x"17",x"12",x"13",x"1b",x"37",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"5b",x"7b",x"5b",x"7b",x"5b",x"3b",x"3b",x"5b",x"5b",x"7b",x"9b",x"bb",x"9b",x"9b",x"9b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"37",x"37",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"12",x"12",x"17",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"32",x"0e",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"12",x"1b",x"13",x"0e",x"12",x"1b",x"17",x"3b",x"17",x"37",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"3b",x"5b",x"3b",x"5b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"0e",x"12",x"1b",x"1b",x"17",x"17",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"12",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"12",x"17",x"1b",x"1b",x"13",x"1b",x"12",x"0e",x"12",x"1b",x"1b",x"1b",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"37",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"5b",x"5b",x"9b",x"9b",x"9b",x"9b",x"5b",x"7b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"0a",x"13",x"1b",x"1b",x"1b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"0e",x"13",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"12",x"12",x"13",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"12",x"0a",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"0e",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"0e",x"0e",x"12",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"13",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"0e",x"0a",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"0e",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"13",x"0e",x"12",x"0e",x"12",x"12",x"12",x"0e",x"32",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"57",x"5b",x"3b",x"5b",x"5b",x"5b",x"3b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"0e",x"12",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"0e",x"0a",x"12",x"12",x"0e",x"12",x"1b",x"3b",x"1b",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"0e",x"37",x"3b",x"3b",x"3b",x"37",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"57",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"12",x"13",x"1b",x"1b",x"1b",x"1b",x"1b",x"12",x"0a",x"12",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"37",x"3b",x"3b",x"3b",x"37",x"12",x"0e",x"37",x"3b",x"3b",x"3b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"13",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"32",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"0e",x"0e",x"17",x"17",x"17",x"1b",x"17",x"0e",x"0a",x"12",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"0e",x"0e",x"0e",x"0e",x"13",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"3b",x"37",x"3b",x"37",x"12",x"0e",x"3b",x"3b",x"3b",x"37",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"13",x"17",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"12",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"3b",x"17",x"17",x"17",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"12",x"12",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"1b",x"17",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"12",x"0e",x"0e",x"0e",x"17",x"1b",x"13",x"0e",x"0a",x"12",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"0e",x"0e",x"0a",x"12",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"17",x"3b",x"37",x"3b",x"37",x"0e",x"0e",x"3b",x"3b",x"3b",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"12",x"12",x"0e",x"12",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"13",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"12",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"5b",x"7b",x"7b",x"7b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"13",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0a",x"12",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0a",x"12",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"3b",x"17",x"0e",x"0e",x"3b",x"3b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"13",x"12",x"13",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"1b",x"17",x"13",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"12",x"12",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"1b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"7b",x"9b",x"bb",x"9b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"0e",x"12",x"3b",x"3b",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"13",x"17",x"17",x"12",x"12",x"17",x"1b",x"1b",x"1b",x"37",x"12",x"1b",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"3b",x"37",x"37",x"37",x"5b",x"9b",x"9b",x"bb",x"9b",x"7b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"1b",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"12",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"17",x"1b",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"0e",x"12",x"3b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"13",x"17",x"17",x"12",x"0e",x"17",x"3b",x"1b",x"1b",x"37",x"12",x"1b",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"5b",x"9b",x"9b",x"bb",x"9b",x"7b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"12",x"1b",x"17",x"17",x"17",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"13",x"0e",x"12",x"1b",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"13",x"17",x"0e",x"12",x"17",x"3b",x"17",x"1b",x"37",x"13",x"17",x"3b",x"3b",x"3b",x"37",x"37",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"5b",x"9b",x"9b",x"9b",x"9b",x"7b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"12",x"1b",x"17",x"17",x"17",x"0e",x"13",x"1b",x"17",x"17",x"1b",x"13",x"17",x"12",x"17",x"17",x"0e",x"0e",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"12",x"0e",x"12",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"12",x"17",x"12",x"12",x"17",x"1b",x"17",x"1b",x"1b",x"37",x"17",x"3b",x"3b",x"3b",x"17",x"12",x"12",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"1b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"7b",x"9b",x"bb",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"12",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"0e",x"17",x"12",x"0e",x"0e",x"0a",x"0e",x"13",x"1b",x"17",x"17",x"17",x"0a",x"12",x"17",x"17",x"12",x"1b",x"13",x"17",x"12",x"17",x"17",x"0a",x"0e",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"17",x"1b",x"17",x"17",x"1b",x"37",x"13",x"3b",x"3b",x"3b",x"37",x"12",x"12",x"12",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"37",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"12",x"0e",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"13",x"12",x"13",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"0e",x"0e",x"1b",x"17",x"13",x"12",x"12",x"0e",x"13",x"1b",x"17",x"1b",x"12",x"0a",x"0e",x"17",x"17",x"0e",x"13",x"13",x"1b",x"12",x"17",x"13",x"0a",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"2e",x"12",x"12",x"17",x"13",x"12",x"12",x"12",x"17",x"3b",x"1b",x"17",x"1b",x"1b",x"12",x"3b",x"3b",x"3b",x"37",x"37",x"12",x"17",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"3b",x"1b",x"1b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"13",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"1b",x"1b",x"1b",x"17",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"13",x"0e",x"0e",x"17",x"1b",x"1b",x"1b",x"17",x"12",x"12",x"17",x"17",x"1b",x"12",x"0e",x"0e",x"17",x"17",x"0e",x"0e",x"12",x"17",x"17",x"17",x"12",x"0a",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"12",x"17",x"3b",x"3b",x"37",x"13",x"12",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"37",x"3b",x"5b",x"3b",x"3b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"3b",x"3b",x"37",x"17",x"1b",x"1b",x"17",x"17",x"17",x"12",x"13",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"12",x"0e",x"0e",x"17",x"12",x"0e",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"13",x"17",x"12",x"0a",x"0e",x"0e",x"12",x"12",x"12",x"0a",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"13",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"13",x"17",x"3b",x"17",x"17",x"12",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"3b",x"7b",x"7b",x"5b",x"3b",x"37",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"5b",x"3b",x"3b",x"1b",x"1b",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"12",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"bb",x"bb",x"7b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"17",x"12",x"12",x"17",x"1b",x"17",x"0e",x"0e",x"0e",x"12",x"1b",x"13",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"3b",x"17",x"12",x"12",x"12",x"37",x"1b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"37",x"5b",x"bb",x"9b",x"7b",x"5b",x"3b",x"1b",x"1b",x"1b",x"17",x"3b",x"9b",x"9b",x"7b",x"5b",x"3b",x"1b",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"12",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"9b",x"7b",x"7b",x"5b",x"5b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"1b",x"17",x"17",x"17",x"1b",x"17",x"12",x"12",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"1b",x"17",x"0e",x"12",x"1b",x"13",x"0e",x"0e",x"0a",x"12",x"1b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"12",x"12",x"12",x"13",x"1b",x"3b",x"37",x"3b",x"3b",x"3b",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"5b",x"9b",x"9b",x"5b",x"5b",x"3b",x"17",x"17",x"17",x"1b",x"5b",x"9b",x"9b",x"7b",x"5b",x"3b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"33",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"13",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"12",x"0e",x"0e",x"0e",x"12",x"17",x"1b",x"1b",x"17",x"12",x"12",x"1b",x"12",x"0e",x"0e",x"0a",x"12",x"1b",x"17",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"0e",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"1b",x"3b",x"3b",x"37",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"5b",x"7b",x"7b",x"5b",x"5b",x"3b",x"17",x"17",x"17",x"1b",x"5b",x"9b",x"9b",x"7b",x"5b",x"5b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"33",x"37",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"13",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"13",x"0e",x"0e",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"0e",x"0e",x"0e",x"0a",x"12",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"0e",x"17",x"17",x"12",x"12",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"1b",x"17",x"17",x"17",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"17",x"37",x"17",x"1b",x"1b",x"1b",x"1b",x"37",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"3b",x"3b",x"3b",x"3b",x"17",x"33",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"37",x"37",x"17",x"17",x"17",x"1b",x"3b",x"5b",x"5b",x"5b",x"57",x"3b",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"3b",x"3b",x"1b",x"1b",x"17",x"1b",x"17",x"1b",x"17",x"12",x"12",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"0e",x"0a",x"0a",x"0e",x"17",x"16",x"13",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"1b",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"0e",x"12",x"12",x"0e",x"0e",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"17",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"37",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"13",x"13",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"13",x"12",x"12",x"12",x"12",x"37",x"1b",x"17",x"17",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"3b",x"5b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"12",x"0e",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"12",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"1b",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"0e",x"12",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"0e",x"12",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"37",x"3b",x"5b",x"5b",x"3b",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"3b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"12",x"13",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"13",x"13",x"37",x"5b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"1b",x"17",x"17",x"17",x"1b",x"13",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"12",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"3b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"37",x"12",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"13",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"37",x"37",x"37",x"1b",x"17",x"17",x"17",x"1b",x"17",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"17",x"13",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"0e",x"0a",x"12",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"32",x"33",x"37",x"17",x"17",x"17",x"1b",x"1b",x"17",x"37",x"37",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"12",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"33",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"33",x"37",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"37",x"3b",x"3b",x"17",x"17",x"37",x"3b",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"5b",x"3b",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"12",x"17",x"13",x"13",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"0e",x"0a",x"12",x"1b",x"17",x"17",x"17",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"13",x"37",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"12",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"37",x"37",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"57",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"37",x"17",x"17",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"5b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"17",x"13",x"13",x"17",x"13",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"12",x"0e",x"0e",x"12",x"1b",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"0e",x"12",x"12",x"0e",x"0e",x"12",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"37",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"17",x"12",x"17",x"1b",x"17",x"37",x"1b",x"17",x"3b",x"37",x"3b",x"37",x"13",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"37",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"3b",x"5b",x"37",x"37",x"5b",x"5b",x"5b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"12",x"12",x"17",x"12",x"0e",x"0e",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"12",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"37",x"37",x"17",x"1b",x"1b",x"17",x"1b",x"17",x"12",x"17",x"1b",x"17",x"17",x"1b",x"37",x"3b",x"3b",x"1b",x"17",x"33",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"37",x"37",x"37",x"37",x"5b",x"37",x"37",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"17",x"17",x"57",x"5b",x"5b",x"37",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"13",x"0a",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0a",x"0e",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"12",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"2e",x"12",x"12",x"32",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"33",x"17",x"1b",x"1b",x"17",x"37",x"37",x"17",x"1b",x"17",x"17",x"1b",x"13",x"12",x"17",x"1b",x"1b",x"17",x"1b",x"37",x"3b",x"3b",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"37",x"37",x"37",x"37",x"5b",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"17",x"57",x"5b",x"57",x"37",x"37",x"37",x"1b",x"1b",x"17",x"17",x"17",x"17",x"0a",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"1b",x"17",x"12",x"0e",x"12",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"0e",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"0a",x"0e",x"13",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"37",x"37",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"12",x"12",x"17",x"1b",x"1b",x"17",x"1b",x"17",x"1b",x"3b",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"37",x"37",x"3b",x"37",x"17",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"bb",x"bb",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"37",x"5b",x"57",x"37",x"37",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"17",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"37",x"37",x"1b",x"12",x"12",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"12",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"37",x"37",x"37",x"17",x"37",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"3b",x"5b",x"57",x"37",x"37",x"3b",x"3b",x"17",x"17",x"17",x"1b",x"17",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"13",x"13",x"12",x"12",x"0e",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"32",x"32",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"32",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"1b",x"1b",x"37",x"37",x"17",x"37",x"12",x"12",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"37",x"12",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"3b",x"17",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"37",x"16",x"3b",x"3b",x"37",x"17",x"17",x"1b",x"17",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0a",x"0e",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"1b",x"1b",x"17",x"37",x"12",x"13",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"7b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"37",x"3b",x"7b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"5b",x"37",x"17",x"37",x"3b",x"3b",x"17",x"17",x"17",x"17",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0a",x"12",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"1b",x"1b",x"37",x"12",x"13",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"13",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"7b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"37",x"5b",x"9b",x"9b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"57",x"57",x"37",x"37",x"17",x"37",x"5b",x"3b",x"3b",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"12",x"0e",x"17",x"12",x"0e",x"0a",x"0e",x"0a",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"13",x"17",x"17",x"12",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"13",x"17",x"17",x"17",x"17",x"13",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"37",x"37",x"37",x"33",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"32",x"12",x"12",x"17",x"17",x"1b",x"17",x"12",x"13",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"13",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"7b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"3b",x"17",x"1b",x"3b",x"5b",x"9b",x"9b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"57",x"37",x"37",x"17",x"37",x"5b",x"3b",x"3b",x"3b",x"17",x"17",x"12",x"0e",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"12",x"0a",x"0e",x"0e",x"0e",x"0a",x"12",x"17",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"12",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"37",x"7b",x"7b",x"37",x"37",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"13",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"13",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"37",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"5b",x"7b",x"9b",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"3b",x"1b",x"17",x"3b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"37",x"37",x"37",x"37",x"37",x"17",x"37",x"5b",x"3b",x"3b",x"3b",x"1b",x"17",x"12",x"0e",x"13",x"17",x"12",x"0e",x"12",x"1b",x"17",x"13",x"12",x"13",x"17",x"17",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"12",x"12",x"13",x"17",x"17",x"12",x"12",x"17",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"57",x"9b",x"9b",x"37",x"37",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"12",x"13",x"17",x"1b",x"17",x"17",x"17",x"3b",x"1b",x"13",x"13",x"1b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"3b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"3b",x"5b",x"5b",x"7b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"17",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"17",x"17",x"37",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"3b",x"3b",x"37",x"37",x"17",x"12",x"0e",x"13",x"17",x"12",x"0e",x"0e",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"17",x"17",x"12",x"12",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"57",x"7b",x"7b",x"37",x"37",x"33",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"1b",x"17",x"3b",x"1b",x"3b",x"1b",x"12",x"17",x"1b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"1b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"37",x"37",x"3b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"37",x"17",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"37",x"17",x"37",x"37",x"17",x"17",x"37",x"37",x"37",x"3b",x"37",x"37",x"5b",x"37",x"37",x"3b",x"12",x"0e",x"13",x"17",x"12",x"0e",x"0e",x"0e",x"17",x"12",x"12",x"17",x"17",x"13",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0a",x"12",x"17",x"12",x"0e",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"32",x"12",x"12",x"32",x"32",x"12",x"12",x"37",x"57",x"37",x"37",x"37",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"12",x"17",x"1b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"3b",x"5b",x"3b",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"17",x"1b",x"17",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"37",x"5b",x"5b",x"37",x"17",x"37",x"37",x"37",x"37",x"37",x"17",x"37",x"5b",x"37",x"3b",x"37",x"16",x"37",x"3b",x"17",x"0e",x"12",x"17",x"12",x"0e",x"0e",x"0e",x"17",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"13",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0a",x"0e",x"12",x"17",x"12",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"37",x"37",x"37",x"37",x"37",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"12",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"37",x"37",x"5b",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"17",x"17",x"1b",x"17",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"37",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"3b",x"37",x"16",x"16",x"37",x"3b",x"17",x"0e",x"12",x"17",x"13",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"0e",x"0a",x"0e",x"0e",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0a",x"0e",x"0e",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"32",x"12",x"12",x"12",x"37",x"37",x"37",x"37",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"1b",x"17",x"1b",x"17",x"12",x"17",x"1b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"37",x"17",x"37",x"3b",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"5b",x"17",x"16",x"37",x"37",x"3b",x"37",x"12",x"12",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"0a",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"33",x"33",x"32",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"37",x"1b",x"1b",x"17",x"12",x"17",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"37",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"3b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"37",x"12",x"37",x"3b",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"17",x"12",x"37",x"3b",x"3b",x"37",x"12",x"12",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"37",x"17",x"1b",x"13",x"12",x"17",x"3b",x"37",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"5b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"5b",x"37",x"37",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"3b",x"3b",x"17",x"12",x"37",x"37",x"37",x"5b",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"17",x"12",x"37",x"3b",x"3b",x"37",x"12",x"12",x"17",x"1b",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"17",x"13",x"13",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"13",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"13",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"1b",x"17",x"12",x"37",x"37",x"37",x"37",x"17",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"17",x"16",x"37",x"3b",x"3b",x"37",x"12",x"12",x"17",x"1b",x"17",x"0e",x"0a",x"0e",x"0a",x"0e",x"13",x"12",x"0a",x"0e",x"0e",x"17",x"17",x"12",x"17",x"13",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"12",x"17",x"17",x"1b",x"1b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"37",x"37",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"12",x"12",x"37",x"17",x"17",x"37",x"5b",x"37",x"37",x"17",x"37",x"37",x"37",x"17",x"17",x"17",x"37",x"3b",x"3b",x"37",x"12",x"12",x"17",x"17",x"17",x"13",x"0e",x"0e",x"12",x"13",x"17",x"12",x"0a",x"0e",x"0e",x"13",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"37",x"17",x"1b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"17",x"37",x"3b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"5b",x"3b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"37",x"37",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"12",x"32",x"16",x"16",x"37",x"5b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"37",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"17",x"12",x"0a",x"0e",x"0e",x"0e",x"17",x"17",x"13",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"32",x"12",x"17",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"3b",x"5b",x"5b",x"3b",x"37",x"57",x"5b",x"3b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"16",x"16",x"32",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"13",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"12",x"12",x"32",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"16",x"17",x"17",x"17",x"37",x"3b",x"3b",x"37",x"37",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"17",x"12",x"0e",x"0e",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"12",x"12",x"12",x"33",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"5b",x"3b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"1b",x"1b",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"37",x"37",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"1b",x"3b",x"1b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"1b",x"17",x"17",x"17",x"17",x"5b",x"5b",x"37",x"3b",x"1b",x"17",x"17",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"37",x"37",x"17",x"37",x"37",x"3b",x"3b",x"37",x"37",x"37",x"12",x"12",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"12",x"0e",x"12",x"17",x"17",x"13",x"12",x"0e",x"0a",x"0e",x"12",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"2e",x"51",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"12",x"12",x"17",x"33",x"33",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"5b",x"5b",x"37",x"5b",x"5b",x"37",x"37",x"37",x"37",x"37",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"13",x"0e",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"12",x"0e",x"13",x"17",x"17",x"17",x"17",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"7b",x"7a",x"7a",x"7a",x"7a",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"1b",x"17",x"17",x"3b",x"7b",x"9b",x"37",x"37",x"1b",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"3b",x"3b",x"37",x"17",x"37",x"12",x"12",x"12",x"17",x"1b",x"17",x"12",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"12",x"0e",x"12",x"17",x"12",x"0e",x"0e",x"0a",x"0a",x"0e",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"2e",x"99",x"51",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"17",x"17",x"32",x"12",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"13",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"13",x"12",x"0e",x"12",x"1b",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"13",x"17",x"17",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"37",x"5b",x"7a",x"9a",x"b9",x"b9",x"b9",x"b9",x"ba",x"9a",x"9a",x"ba",x"9a",x"9a",x"9a",x"9a",x"9a",x"5b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"57",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"17",x"17",x"17",x"17",x"5b",x"9b",x"9b",x"57",x"37",x"3b",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"37",x"16",x"37",x"12",x"12",x"12",x"12",x"17",x"17",x"12",x"1b",x"17",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"2e",x"b9",x"95",x"2e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"2e",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"12",x"33",x"37",x"13",x"12",x"12",x"12",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"5b",x"3b",x"37",x"37",x"37",x"3b",x"5b",x"5b",x"37",x"5b",x"5b",x"3b",x"17",x"12",x"12",x"13",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"13",x"12",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"5b",x"7a",x"9a",x"9a",x"9a",x"9a",x"9a",x"7a",x"7a",x"7a",x"7a",x"7a",x"7a",x"7a",x"7a",x"7a",x"7a",x"7a",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"9b",x"9b",x"7b",x"7b",x"9b",x"7b",x"7b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"12",x"17",x"17",x"37",x"5b",x"9b",x"9b",x"57",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"37",x"37",x"3b",x"37",x"17",x"17",x"37",x"12",x"12",x"12",x"12",x"17",x"17",x"12",x"17",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0a",x"12",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"b9",x"b9",x"71",x"2e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"71",x"75",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"32",x"12",x"33",x"33",x"12",x"17",x"37",x"17",x"33",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"37",x"3b",x"37",x"3b",x"5b",x"3b",x"37",x"3b",x"3b",x"17",x"12",x"0e",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"12",x"12",x"0e",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"7a",x"ba",x"b9",x"b9",x"9a",x"7a",x"37",x"3b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"9b",x"7b",x"9b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"3b",x"37",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"17",x"17",x"17",x"5b",x"7b",x"7b",x"37",x"37",x"17",x"17",x"12",x"12",x"12",x"17",x"37",x"3b",x"3b",x"37",x"37",x"16",x"37",x"3b",x"3b",x"37",x"37",x"37",x"12",x"17",x"37",x"12",x"12",x"12",x"12",x"17",x"17",x"12",x"12",x"12",x"0e",x"12",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"99",x"b8",x"98",x"51",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"95",x"d9",x"b8",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"32",x"33",x"32",x"33",x"17",x"17",x"37",x"37",x"37",x"17",x"17",x"17",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"5b",x"3b",x"37",x"37",x"3b",x"5b",x"37",x"17",x"17",x"17",x"1b",x"17",x"12",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"7a",x"ba",x"b9",x"9a",x"7a",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"37",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"17",x"17",x"17",x"3b",x"5b",x"5b",x"3b",x"37",x"33",x"12",x"12",x"12",x"17",x"17",x"17",x"37",x"3b",x"3b",x"37",x"16",x"17",x"37",x"3b",x"37",x"17",x"17",x"16",x"17",x"37",x"12",x"12",x"12",x"12",x"13",x"17",x"12",x"32",x"12",x"0e",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0a",x"0e",x"12",x"17",x"13",x"17",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"99",x"99",x"98",x"99",x"51",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"52",x"b9",x"b9",x"94",x"95",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"33",x"32",x"33",x"32",x"33",x"17",x"17",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"37",x"3b",x"3b",x"17",x"12",x"17",x"17",x"1b",x"17",x"12",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"13",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"1b",x"17",x"3b",x"5a",x"9a",x"b9",x"9a",x"5a",x"37",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"37",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"37",x"32",x"12",x"13",x"17",x"17",x"1b",x"17",x"17",x"1b",x"3b",x"37",x"17",x"16",x"17",x"37",x"37",x"17",x"17",x"16",x"17",x"37",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"13",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"99",x"95",x"95",x"98",x"99",x"51",x"2e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"32",x"95",x"b9",x"b8",x"74",x"75",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"33",x"32",x"32",x"33",x"33",x"13",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"3b",x"3b",x"37",x"37",x"37",x"12",x"12",x"17",x"17",x"1b",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"13",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"37",x"1b",x"37",x"7a",x"b9",x"b9",x"9a",x"3b",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"37",x"37",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0a",x"13",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"3b",x"37",x"12",x"16",x"17",x"37",x"37",x"17",x"17",x"17",x"37",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"17",x"17",x"17",x"13",x"17",x"17",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"95",x"95",x"95",x"98",x"98",x"98",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"2e",x"95",x"b9",x"99",x"94",x"74",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"33",x"33",x"33",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"37",x"37",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"3b",x"37",x"37",x"12",x"12",x"12",x"17",x"17",x"1b",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"13",x"17",x"17",x"17",x"13",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"1b",x"37",x"7a",x"b9",x"b9",x"7a",x"3b",x"37",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"37",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0a",x"13",x"17",x"17",x"17",x"13",x"0e",x"17",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"17",x"17",x"17",x"17",x"17",x"16",x"17",x"37",x"3b",x"37",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0a",x"75",x"b9",x"95",x"74",x"b8",x"98",x"99",x"51",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0a",x"75",x"99",x"98",x"74",x"74",x"98",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"33",x"33",x"33",x"33",x"33",x"37",x"37",x"17",x"17",x"37",x"37",x"37",x"17",x"17",x"37",x"37",x"37",x"37",x"3b",x"37",x"37",x"37",x"3b",x"37",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"13",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"1b",x"3b",x"7a",x"b9",x"b9",x"7a",x"3b",x"17",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"9b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"13",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"3b",x"1b",x"17",x"0e",x"12",x"17",x"17",x"17",x"12",x"0e",x"13",x"13",x"12",x"17",x"13",x"12",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"16",x"16",x"17",x"37",x"3b",x"3b",x"37",x"12",x"12",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0a",x"51",x"b9",x"95",x"71",x"95",x"98",x"98",x"99",x"51",x"0e",x"0a",x"0e",x"0e",x"0a",x"32",x"99",x"98",x"98",x"74",x"74",x"99",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"33",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"37",x"37",x"37",x"37",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"17",x"17",x"17",x"12",x"0e",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"1b",x"17",x"5b",x"b9",x"b9",x"7a",x"3b",x"1b",x"37",x"3b",x"3b",x"1b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"12",x"17",x"17",x"17",x"17",x"5b",x"9b",x"9b",x"7b",x"5b",x"1b",x"17",x"0e",x"0e",x"17",x"17",x"17",x"12",x"0e",x"12",x"13",x"12",x"13",x"0e",x"0e",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"16",x"17",x"37",x"37",x"37",x"37",x"37",x"12",x"12",x"17",x"17",x"12",x"13",x"17",x"12",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"2e",x"99",x"b9",x"75",x"71",x"b9",x"99",x"98",x"98",x"51",x"0a",x"0e",x"0e",x"0a",x"95",x"99",x"78",x"78",x"74",x"74",x"75",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"33",x"33",x"33",x"37",x"37",x"37",x"37",x"17",x"17",x"37",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"13",x"12",x"0e",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"13",x"0e",x"17",x"17",x"17",x"12",x"0e",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"5b",x"9a",x"b9",x"7a",x"3b",x"17",x"1b",x"1b",x"3b",x"17",x"37",x"3b",x"3b",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"3b",x"5b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"12",x"17",x"17",x"17",x"17",x"7b",x"9b",x"9b",x"9b",x"5b",x"1b",x"3b",x"32",x"0e",x"13",x"17",x"17",x"13",x"0e",x"0e",x"13",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"37",x"37",x"37",x"17",x"16",x"17",x"17",x"17",x"37",x"17",x"12",x"16",x"17",x"17",x"13",x"17",x"17",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"95",x"dd",x"95",x"50",x"99",x"99",x"98",x"98",x"75",x"31",x"0a",x"0a",x"2e",x"99",x"75",x"75",x"75",x"75",x"75",x"55",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"13",x"13",x"33",x"33",x"37",x"37",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"12",x"12",x"0e",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"0e",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"9a",x"b9",x"9a",x"3b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"37",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"37",x"1b",x"3b",x"3b",x"3b",x"37",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"37",x"5b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"13",x"17",x"17",x"17",x"7b",x"7b",x"7b",x"9b",x"5b",x"17",x"3b",x"32",x"0e",x"13",x"17",x"17",x"13",x"0e",x"0e",x"12",x"0e",x"0a",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"12",x"16",x"16",x"12",x"17",x"17",x"17",x"16",x"17",x"17",x"13",x"13",x"17",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"13",x"0e",x"13",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"13",x"12",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"75",x"bd",x"99",x"70",x"74",x"99",x"95",x"79",x"98",x"75",x"2e",x"0a",x"71",x"94",x"74",x"75",x"75",x"75",x"51",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"33",x"33",x"33",x"37",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"13",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"0e",x"13",x"17",x"12",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"5a",x"b9",x"b9",x"5b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"12",x"17",x"17",x"1b",x"7b",x"9b",x"7b",x"7b",x"5b",x"1b",x"1b",x"32",x"0e",x"13",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"17",x"16",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"33",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"51",x"99",x"b9",x"95",x"4c",x"99",x"95",x"74",x"74",x"74",x"51",x"2e",x"95",x"75",x"74",x"75",x"75",x"50",x"51",x"2d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"33",x"33",x"33",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"32",x"33",x"33",x"13",x"13",x"33",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"17",x"13",x"17",x"17",x"17",x"13",x"12",x"17",x"12",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"5b",x"9a",x"b9",x"7a",x"1b",x"17",x"17",x"17",x"37",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"37",x"37",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"37",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"12",x"17",x"17",x"1b",x"3b",x"5b",x"7b",x"5b",x"3b",x"1b",x"1b",x"37",x"0e",x"13",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"13",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"12",x"12",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"2e",x"75",x"b9",x"99",x"50",x"75",x"99",x"75",x"75",x"75",x"55",x"51",x"75",x"75",x"75",x"74",x"50",x"50",x"51",x"2e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"33",x"33",x"37",x"37",x"37",x"37",x"37",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"17",x"17",x"0e",x"13",x"12",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"7a",x"b9",x"9a",x"3b",x"1b",x"17",x"17",x"17",x"37",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"37",x"37",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"37",x"17",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"5b",x"5b",x"3b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"5b",x"3b",x"5b",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"12",x"17",x"17",x"1b",x"1b",x"3b",x"5b",x"3b",x"17",x"1b",x"1b",x"17",x"0e",x"12",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"17",x"17",x"17",x"16",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"17",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"51",x"b8",x"99",x"95",x"50",x"75",x"75",x"75",x"75",x"75",x"74",x"74",x"75",x"55",x"50",x"4c",x"50",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"36",x"36",x"36",x"36",x"37",x"37",x"37",x"37",x"37",x"37",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"13",x"0e",x"0e",x"12",x"13",x"17",x"17",x"17",x"13",x"17",x"17",x"13",x"12",x"12",x"0e",x"12",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"37",x"37",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"5a",x"b9",x"b9",x"7b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"37",x"37",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"13",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0a",x"0a",x"0a",x"0a",x"0a",x"0a",x"0a",x"0a",x"0e",x"0e",x"0a",x"51",x"99",x"99",x"99",x"50",x"75",x"75",x"75",x"54",x"74",x"75",x"54",x"75",x"50",x"51",x"4d",x"4c",x"51",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"32",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"37",x"37",x"37",x"37",x"37",x"37",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"0e",x"17",x"17",x"13",x"0e",x"12",x"12",x"12",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"17",x"17",x"17",x"13",x"13",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"9a",x"b9",x"9a",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"3b",x"37",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"17",x"37",x"5b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"13",x"17",x"17",x"3b",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"12",x"0e",x"12",x"17",x"12",x"0e",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"17",x"17",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"35",x"75",x"98",x"99",x"74",x"50",x"75",x"75",x"55",x"75",x"55",x"55",x"51",x"50",x"50",x"4c",x"4c",x"51",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"32",x"32",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"5a",x"3a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"36",x"57",x"57",x"57",x"36",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"13",x"12",x"33",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"3b",x"3b",x"17",x"17",x"37",x"37",x"37",x"17",x"37",x"17",x"1b",x"37",x"13",x"12",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"7a",x"b9",x"b9",x"5a",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"3b",x"37",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"3b",x"37",x"3b",x"3b",x"3b",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"3b",x"37",x"3b",x"17",x"1b",x"1b",x"0e",x"0e",x"12",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"15",x"15",x"15",x"15",x"16",x"15",x"16",x"16",x"15",x"55",x"74",x"75",x"75",x"31",x"51",x"75",x"75",x"55",x"51",x"55",x"50",x"51",x"50",x"4c",x"4c",x"51",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"0e",x"0e",x"0e",x"0e"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"3a",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"36",x"36",x"36",x"36",x"36",x"36",x"56",x"56",x"56",x"56",x"56",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"37",x"37",x"37",x"37",x"17",x"17",x"37",x"37",x"3b",x"3b",x"37",x"17",x"1b",x"3b",x"17",x"37",x"37",x"37",x"37",x"17",x"1b",x"1b",x"17",x"1b",x"17",x"12",x"13",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"37",x"9a",x"b9",x"9a",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"17",x"3b",x"3b",x"1b",x"1b",x"17",x"0e",x"0e",x"0e",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"16",x"16",x"16",x"16",x"16",x"15",x"16",x"16",x"35",x"71",x"74",x"75",x"75",x"2c",x"50",x"75",x"51",x"51",x"51",x"50",x"4c",x"51",x"2c",x"2c",x"31",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"3a",x"3a",x"3a",x"3a",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"16",x"36",x"5a",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5a",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"37",x"37",x"1b",x"3b",x"37",x"1b",x"3b",x"1b",x"37",x"37",x"37",x"37",x"37",x"17",x"17",x"1b",x"17",x"1b",x"17",x"13",x"13",x"17",x"13",x"17",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"5b",x"b9",x"b9",x"5a",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"5b",x"3b",x"3b",x"3b",x"37",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"33",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"11",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"35",x"70",x"75",x"75",x"50",x"50",x"51",x"55",x"51",x"51",x"4c",x"4c",x"51",x"4c",x"2c",x"31",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"36",x"36",x"36",x"36",x"36",x"16",x"16",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"3a",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"5a",x"56",x"56",x"5a",x"5a",x"5a",x"5a",x"5a",x"5b",x"5b",x"5a",x"5a",x"5a",x"5a",x"5a",x"56",x"56",x"36",x"37",x"1b",x"1b",x"1b",x"1b",x"3b",x"17",x"37",x"37",x"37",x"17",x"13",x"17",x"17",x"17",x"17",x"1b",x"17",x"37",x"13",x"17",x"13",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"9a",x"b9",x"9a",x"37",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"37",x"3b",x"3b",x"3b",x"37",x"37",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"17",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"16",x"1a",x"16",x"16",x"1a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"16",x"16",x"16",x"15",x"15",x"16",x"16",x"16",x"16",x"15",x"51",x"50",x"75",x"51",x"50",x"50",x"51",x"50",x"4c",x"4c",x"2c",x"4c",x"2c",x"2c",x"31",x"16",x"16",x"16",x"15",x"16",x"16",x"16",x"16",x"16",x"35",x"16",x"16",x"16",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"16",x"36",x"36",x"36",x"16",x"16",x"16",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"5a",x"5a",x"5a",x"56",x"5a",x"5a",x"5a",x"5a",x"56",x"56",x"37",x"3b",x"1b",x"17",x"1b",x"1b",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"57",x"b9",x"b9",x"5a",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"16",x"16",x"15",x"16",x"16",x"16",x"16",x"16",x"15",x"11",x"11",x"50",x"50",x"50",x"50",x"2c",x"4c",x"50",x"4c",x"2c",x"2c",x"2c",x"2c",x"2c",x"31",x"12",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"16",x"75",x"16",x"16",x"16",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"15",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"16",x"36",x"36",x"16",x"16",x"16",x"16",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"5a",x"56",x"56",x"5a",x"5a",x"5a",x"5a",x"3b",x"3b",x"17",x"17",x"17",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"13",x"37",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"12",x"13",x"17",x"17",x"17",x"37",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"7a",x"b9",x"b9",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"1b",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"13",x"17",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"16",x"16",x"15",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"16",x"15",x"11",x"12",x"16",x"15",x"16",x"12",x"11",x"11",x"11",x"31",x"51",x"50",x"4c",x"2c",x"2c",x"4c",x"4d",x"2c",x"2d",x"28",x"28",x"2d",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"16",x"94",x"35",x"16",x"16",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"15",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"12",x"16",x"16",x"12",x"11",x"12",x"16",x"16",x"12",x"11",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"37",x"37",x"37",x"36",x"36",x"16",x"16",x"36",x"3b",x"5b",x"56",x"56",x"5a",x"5a",x"5a",x"5a",x"5a",x"3b",x"37",x"17",x"17",x"32",x"37",x"37",x"37",x"17",x"37",x"37",x"33",x"37",x"37",x"17",x"1b",x"17",x"37",x"37",x"1b",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"99",x"b9",x"7a",x"37",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"5b",x"9b",x"37",x"17",x"1b",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"3b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"17",x"37",x"3b",x"3b",x"37",x"37",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"1a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"16",x"12",x"12",x"12",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"16",x"31",x"4d",x"50",x"4c",x"2c",x"2c",x"4c",x"2c",x"2d",x"28",x"2c",x"31",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"35",x"94",x"55",x"16",x"16",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0a",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"12",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"16",x"36",x"37",x"36",x"36",x"36",x"16",x"17",x"37",x"36",x"5a",x"5a",x"5a",x"5a",x"5a",x"56",x"56",x"56",x"5a",x"5a",x"37",x"37",x"17",x"36",x"37",x"33",x"33",x"17",x"37",x"33",x"37",x"17",x"37",x"17",x"17",x"17",x"37",x"33",x"17",x"17",x"37",x"17",x"17",x"17",x"37",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"5b",x"b9",x"b9",x"57",x"17",x"17",x"17",x"37",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"da",x"f9",x"7b",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"13",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"31",x"4c",x"4c",x"28",x"2c",x"2c",x"2d",x"2c",x"2d",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"55",x"94",x"75",x"16",x"16",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"15",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"5a",x"5a",x"5a",x"5a",x"5a",x"56",x"56",x"5a",x"56",x"56",x"5a",x"3b",x"17",x"17",x"17",x"33",x"33",x"17",x"33",x"33",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"33",x"17",x"17",x"37",x"37",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"17",x"17",x"7a",x"b9",x"99",x"37",x"17",x"17",x"17",x"37",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"f9",x"f9",x"ba",x"37",x"17",x"1b",x"1b",x"1b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"13",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"1b",x"1b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"7b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"13",x"12",x"12",x"12",x"12",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"1a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"16",x"16",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"31",x"2d",x"2d",x"28",x"2c",x"28",x"2d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"75",x"74",x"75",x"35",x"12",x"12",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"56",x"5a",x"5a",x"5a",x"5a",x"56",x"56",x"56",x"36",x"5a",x"5a",x"56",x"56",x"5a",x"3b",x"37",x"17",x"17",x"33",x"33",x"17",x"33",x"33",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"37",x"33",x"33",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"33",x"13",x"12",x"32",x"17",x"37",x"ba",x"b9",x"7a",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"f9",x"f9",x"f9",x"7b",x"17",x"1b",x"1b",x"17",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"13",x"17",x"17",x"12",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"1b",x"3b",x"3b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"5b",x"7b",x"7b",x"7b",x"5b",x"37",x"37",x"3b",x"3b",x"3b",x"37",x"5b",x"3b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"13",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"16",x"16",x"16",x"12",x"11",x"15",x"16",x"16",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"31",x"2d",x"28",x"28",x"11",x"16",x"11",x"11",x"11",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"75",x"70",x"74",x"31",x"12",x"11",x"11",x"12"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0a",x"0a",x"0e",x"0e",x"12",x"12",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"56",x"56",x"5a",x"56",x"56",x"5a",x"5a",x"5a",x"56",x"5a",x"5a",x"36",x"5b",x"5a",x"56",x"5a",x"3a",x"37",x"17",x"17",x"37",x"33",x"33",x"33",x"33",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"32",x"17",x"17",x"33",x"32",x"13",x"17",x"37",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"12",x"33",x"13",x"12",x"17",x"17",x"5b",x"b9",x"b9",x"57",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"57",x"f9",x"d9",x"f9",x"9a",x"37",x"1b",x"17",x"17",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"13",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"3b",x"3b",x"37",x"3b",x"37",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"12",x"11",x"11",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"15",x"15",x"16",x"11",x"08",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"31",x"70",x"50",x"74",x"31",x"12",x"11",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"15",x"15",x"15",x"11",x"11",x"11",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"16",x"16",x"16",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"56",x"56",x"5a",x"5a",x"5a",x"56",x"5a",x"5a",x"56",x"56",x"5a",x"5a",x"36",x"57",x"5a",x"56",x"5a",x"5a",x"56",x"37",x"17",x"17",x"13",x"33",x"33",x"13",x"33",x"37",x"17",x"17",x"17",x"17",x"17",x"32",x"17",x"17",x"33",x"32",x"12",x"33",x"33",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"12",x"12",x"33",x"12",x"17",x"17",x"37",x"7a",x"b9",x"b9",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"77",x"f9",x"b5",x"f9",x"da",x"5b",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"5b",x"3b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"3b",x"3b",x"3b",x"3b",x"37",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"56",x"57",x"32",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"36",x"36",x"1a",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"16",x"16",x"16",x"16",x"0c",x"0d",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"55",x"50",x"2c",x"74",x"35",x"12",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"15",x"15",x"15",x"16",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"16",x"16",x"16",x"15",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"3a",x"5a",x"5a",x"56",x"5a",x"56",x"56",x"56",x"56",x"56",x"5a",x"36",x"5a",x"56",x"56",x"56",x"56",x"56",x"5a",x"37",x"17",x"17",x"17",x"33",x"33",x"17",x"32",x"33",x"17",x"17",x"37",x"17",x"17",x"16",x"17",x"1b",x"37",x"32",x"13",x"13",x"33",x"13",x"13",x"17",x"33",x"37",x"37",x"33",x"32",x"12",x"33",x"12",x"17",x"17",x"37",x"99",x"b9",x"9a",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"9a",x"f9",x"b5",x"f9",x"f9",x"7a",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"1b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"3b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"3b",x"3b",x"3b",x"3b",x"17",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"32",x"9b",x"7b",x"37",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"36",x"3a",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"16",x"0d",x"0d",x"11",x"12",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"75",x"2c",x"2c",x"74",x"55",x"16",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"15",x"15",x"15",x"16",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"56",x"56",x"56",x"56",x"5a",x"5a",x"36",x"56",x"5a",x"56",x"5a",x"37",x"17",x"37",x"33",x"33",x"33",x"12",x"12",x"33",x"33",x"17",x"37",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"13",x"12",x"33",x"13",x"33",x"17",x"17",x"17",x"17",x"12",x"32",x"12",x"32",x"17",x"17",x"17",x"56",x"b9",x"b9",x"7a",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"fa",x"f9",x"b5",x"f9",x"f9",x"ba",x"3b",x"1b",x"1b",x"1b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"37",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"12",x"37",x"17",x"1b",x"17",x"17",x"37",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"37",x"17",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"57",x"3b",x"3b",x"37",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"12",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"57",x"9b",x"9b",x"37",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"0d",x"0c",x"0d",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"70",x"2c",x"2c",x"70",x"55",x"11",x"12",x"12",x"12"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"15",x"15",x"16",x"16",x"16",x"16",x"11",x"11",x"12",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"56",x"5a",x"36",x"36",x"56",x"36",x"5a",x"37",x"32",x"33",x"33",x"33",x"33",x"12",x"17",x"33",x"33",x"17",x"17",x"17",x"17",x"17",x"12",x"37",x"17",x"17",x"17",x"12",x"32",x"13",x"33",x"17",x"13",x"12",x"12",x"12",x"32",x"12",x"33",x"17",x"17",x"17",x"5a",x"b9",x"b9",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"7a",x"f9",x"f9",x"b5",x"d9",x"f9",x"fa",x"7b",x"17",x"1b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"37",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"17",x"37",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"37",x"3b",x"3b",x"3b",x"37",x"17",x"37",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"37",x"3b",x"3b",x"37",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"37",x"77",x"77",x"37",x"37",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"16",x"3a",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"0c",x"0d",x"12",x"11",x"12",x"11",x"11",x"11",x"11",x"31",x"51",x"50",x"2c",x"2c",x"50",x"51",x"31",x"12",x"11",x"11"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0e",x"0e",x"12",x"11",x"16",x"16",x"16",x"15",x"11",x"11",x"12",x"16",x"16",x"16",x"11",x"0d",x"11",x"16",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"56",x"3a",x"36",x"36",x"56",x"5a",x"36",x"12",x"33",x"33",x"33",x"33",x"13",x"17",x"13",x"33",x"17",x"17",x"17",x"17",x"17",x"32",x"17",x"17",x"17",x"17",x"12",x"12",x"33",x"33",x"13",x"12",x"32",x"33",x"33",x"33",x"12",x"17",x"17",x"17",x"37",x"7a",x"b9",x"99",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"57",x"da",x"f9",x"f9",x"b5",x"d9",x"f9",x"f9",x"ba",x"17",x"17",x"3b",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"17",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"37",x"3b",x"3b",x"3b",x"37",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"3b",x"3b",x"37",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"37",x"36",x"33",x"37",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"1a",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"11",x"12",x"12",x"11",x"11",x"0d",x"11",x"11",x"0c",x"0d",x"12",x"12",x"12",x"11",x"11",x"11",x"12",x"31",x"50",x"2c",x"0c",x"2c",x"50",x"51",x"31",x"11",x"11",x"11"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0e",x"0e",x"12",x"12",x"11",x"16",x"15",x"15",x"15",x"15",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"56",x"56",x"36",x"36",x"36",x"5a",x"36",x"36",x"12",x"33",x"33",x"33",x"33",x"33",x"13",x"13",x"33",x"17",x"17",x"17",x"37",x"17",x"33",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"12",x"32",x"32",x"33",x"12",x"13",x"17",x"17",x"17",x"17",x"57",x"9a",x"b9",x"7a",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"76",x"f9",x"f9",x"f9",x"b5",x"d9",x"f9",x"f9",x"da",x"37",x"1b",x"1b",x"3b",x"37",x"3b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"37",x"37",x"17",x"3b",x"1b",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"17",x"17",x"37",x"3b",x"3b",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"17",x"37",x"37",x"37",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"37",x"17",x"37",x"33",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"36",x"16",x"16",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"55",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"0d",x"0d",x"11",x"11",x"11",x"11",x"0d",x"11",x"0c",x"0d",x"12",x"11",x"11",x"11",x"12",x"11",x"31",x"51",x"50",x"2c",x"08",x"2c",x"50",x"51",x"31",x"11",x"11",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"15",x"16",x"16",x"15",x"15",x"15",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"5a",x"36",x"36",x"36",x"3a",x"36",x"36",x"12",x"12",x"33",x"33",x"33",x"33",x"32",x"13",x"13",x"33",x"17",x"17",x"17",x"37",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"32",x"33",x"33",x"13",x"17",x"17",x"17",x"17",x"17",x"56",x"b9",x"99",x"56",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"37",x"96",x"f9",x"f9",x"f9",x"b5",x"d9",x"f9",x"fd",x"da",x"5b",x"1b",x"1b",x"3b",x"37",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"12",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"17",x"17",x"37",x"3b",x"37",x"17",x"17",x"37",x"3b",x"37",x"3b",x"3b",x"37",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"37",x"37",x"17",x"17",x"17",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"33",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"1a",x"1a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"b9",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"0d",x"0d",x"11",x"11",x"11",x"12",x"0d",x"11",x"08",x"0d",x"11",x"11",x"11",x"11",x"11",x"12",x"31",x"51",x"2c",x"2c",x"08",x"2d",x"50",x"51",x"31",x"11",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"12",x"12",x"16",x"11",x"12",x"16",x"16",x"15",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"56",x"5a",x"56",x"56",x"56",x"56",x"5a",x"56",x"56",x"36",x"36",x"3a",x"5a",x"3a",x"36",x"12",x"12",x"12",x"33",x"33",x"33",x"33",x"32",x"12",x"12",x"33",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"33",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"76",x"b8",x"99",x"56",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"13",x"13",x"13",x"56",x"b5",x"f8",x"f9",x"fd",x"b5",x"da",x"fe",x"fe",x"da",x"7b",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"13",x"17",x"13",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"17",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"3b",x"37",x"17",x"17",x"3b",x"3b",x"37",x"3b",x"37",x"5b",x"5b",x"5b",x"3b",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"35",x"d9",x"75",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"0d",x"08",x"0d",x"11",x"11",x"11",x"11",x"11",x"12",x"31",x"4c",x"2d",x"28",x"08",x"2c",x"50",x"51",x"35",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"11",x"16",x"16",x"16",x"16",x"11",x"15",x"15",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"56",x"5a",x"56",x"56",x"56",x"56",x"56",x"36",x"56",x"36",x"3a",x"5a",x"36",x"36",x"12",x"12",x"12",x"12",x"13",x"33",x"33",x"33",x"33",x"32",x"32",x"33",x"17",x"17",x"17",x"17",x"17",x"33",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"33",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"75",x"b8",x"75",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"13",x"13",x"13",x"56",x"d5",x"f8",x"f9",x"f9",x"b5",x"da",x"fe",x"fd",x"da",x"57",x"1b",x"17",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"12",x"0e",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"1b",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"37",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"5b",x"3b",x"37",x"17",x"1b",x"17",x"17",x"3b",x"3b",x"37",x"37",x"17",x"3b",x"37",x"17",x"17",x"37",x"37",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"57",x"57",x"33",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"55",x"d9",x"99",x"55",x"35",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"0d",x"08",x"0d",x"11",x"12",x"12",x"15",x"16",x"31",x"2c",x"2c",x"2c",x"28",x"0c",x"2c",x"50",x"51",x"15",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"15",x"15",x"15",x"11",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"11",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"56",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"13",x"33",x"33",x"33",x"33",x"32",x"32",x"33",x"13",x"17",x"17",x"17",x"17",x"33",x"32",x"32",x"17",x"17",x"17",x"17",x"17",x"17",x"33",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"36",x"95",x"b8",x"75",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"36",x"b5",x"f8",x"f8",x"f8",x"b5",x"d9",x"f9",x"fd",x"da",x"57",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"37",x"37",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"13",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"17",x"1b",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"3b",x"17",x"37",x"3b",x"3b",x"3b",x"37",x"17",x"3b",x"37",x"17",x"17",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"13",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"7b",x"9b",x"37",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"1a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"75",x"b9",x"b9",x"99",x"75",x"55",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"0d",x"08",x"0c",x"11",x"16",x"16",x"16",x"16",x"31",x"2c",x"2c",x"2c",x"28",x"0c",x"2c",x"70",x"51",x"11",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0a",x"0e",x"0e",x"12",x"12",x"11",x"11",x"11",x"15",x"16",x"16",x"16",x"15",x"11",x"12",x"16",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"36",x"16",x"36",x"36",x"36",x"36",x"3a",x"36",x"36",x"36",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"3a",x"36",x"36",x"3a",x"5a",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"33",x"33",x"33",x"32",x"32",x"33",x"13",x"32",x"33",x"17",x"17",x"33",x"32",x"12",x"33",x"17",x"17",x"37",x"17",x"1b",x"33",x"17",x"17",x"13",x"13",x"13",x"13",x"12",x"13",x"56",x"99",x"98",x"75",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"33",x"95",x"d4",x"d4",x"d4",x"b4",x"d4",x"d9",x"fa",x"ba",x"57",x"17",x"1b",x"1b",x"1b",x"1b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"5b",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"33",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"5b",x"5b",x"5b",x"5b",x"3b",x"1b",x"37",x"1b",x"37",x"17",x"3b",x"37",x"37",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"17",x"17",x"17",x"3b",x"5b",x"37",x"37",x"3b",x"5b",x"3b",x"37",x"17",x"3b",x"37",x"17",x"37",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"37",x"9b",x"9b",x"57",x"37",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"99",x"95",x"b9",x"99",x"99",x"99",x"99",x"75",x"75",x"55",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"08",x"08",x"11",x"16",x"16",x"16",x"31",x"2c",x"2c",x"2c",x"28",x"08",x"2c",x"2c",x"70",x"51",x"15",x"16",x"16",x"15"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"15",x"15",x"15",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"16",x"12",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"36",x"36",x"36",x"3a",x"3a",x"36",x"36",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"5a",x"5a",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"33",x"33",x"13",x"32",x"32",x"32",x"33",x"33",x"33",x"33",x"17",x"17",x"33",x"33",x"12",x"32",x"17",x"17",x"37",x"17",x"17",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"13",x"55",x"98",x"99",x"56",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"76",x"d4",x"d4",x"d4",x"b4",x"d4",x"d4",x"d5",x"ba",x"37",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"37",x"17",x"17",x"37",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"37",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"37",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"5b",x"5b",x"3b",x"17",x"1b",x"1b",x"3b",x"17",x"17",x"1b",x"37",x"37",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"37",x"3b",x"37",x"17",x"17",x"3b",x"3b",x"5b",x"37",x"37",x"3b",x"5b",x"3b",x"37",x"17",x"37",x"17",x"17",x"37",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"37",x"57",x"57",x"37",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"99",x"95",x"95",x"b9",x"b9",x"99",x"99",x"99",x"99",x"75",x"55",x"55",x"35",x"32",x"12",x"12",x"12",x"12",x"12",x"0d",x"0c",x"11",x"16",x"12",x"16",x"31",x"2c",x"2c",x"28",x"28",x"08",x"2c",x"2c",x"70",x"31",x"16",x"16",x"12",x"0d"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"11",x"15",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"56",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"36",x"36",x"36",x"3a",x"3a",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"33",x"33",x"13",x"33",x"32",x"12",x"33",x"33",x"33",x"33",x"33",x"37",x"33",x"33",x"33",x"33",x"17",x"17",x"17",x"13",x"12",x"0e",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"13",x"75",x"98",x"99",x"56",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"36",x"b5",x"d4",x"d4",x"b4",x"b4",x"d4",x"d5",x"76",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"37",x"37",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"37",x"37",x"37",x"37",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"37",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"37",x"1b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"5b",x"37",x"37",x"37",x"5b",x"3b",x"37",x"17",x"37",x"17",x"37",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"36",x"37",x"12",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"95",x"99",x"95",x"b9",x"b9",x"99",x"99",x"99",x"99",x"99",x"98",x"99",x"75",x"55",x"31",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"12",x"12",x"11",x"2c",x"2c",x"2c",x"28",x"2c",x"08",x"2c",x"4d",x"50",x"31",x"16",x"12",x"0d",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"15",x"12",x"12",x"15",x"15",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"11",x"0d",x"0d",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"0d",x"0d",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"36",x"3a",x"5a",x"5a",x"3a",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"33",x"33",x"13",x"33",x"32",x"12",x"33",x"33",x"13",x"13",x"32",x"12",x"33",x"13",x"33",x"13",x"12",x"12",x"13",x"12",x"0e",x"12",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"33",x"79",x"98",x"75",x"32",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"56",x"d4",x"d4",x"b4",x"d4",x"d4",x"96",x"37",x"17",x"1b",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"1b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"37",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"37",x"33",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"37",x"37",x"12",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"37",x"17",x"3b",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"37",x"5b",x"3b",x"37",x"37",x"37",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"37",x"37",x"33",x"37",x"12",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"75",x"b9",x"75",x"99",x"b9",x"99",x"99",x"99",x"75",x"79",x"79",x"75",x"75",x"75",x"75",x"55",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"12",x"12",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"2c",x"2c",x"51",x"50",x"31",x"11",x"0d",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"11",x"15",x"15",x"12",x"12",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"11",x"0d",x"0d",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"0d",x"0d",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"3a",x"3a",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"3a",x"36",x"36",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"33",x"33",x"33",x"33",x"33",x"12",x"32",x"33",x"33",x"33",x"33",x"32",x"33",x"13",x"12",x"12",x"0e",x"0e",x"13",x"12",x"0e",x"12",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"32",x"79",x"98",x"75",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"95",x"d4",x"b4",x"d4",x"95",x"36",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"33",x"17",x"37",x"33",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"17",x"17",x"17",x"13",x"13",x"12",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"37",x"37",x"12",x"12",x"17",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"37",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"37",x"5b",x"3b",x"37",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0a",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"35",x"b9",x"95",x"95",x"99",x"b9",x"99",x"79",x"75",x"75",x"75",x"75",x"75",x"74",x"75",x"75",x"55",x"31",x"12",x"0d",x"0d",x"0d",x"16",x"11",x"2d",x"2d",x"2d",x"2d",x"2d",x"0c",x"2c",x"2c",x"51",x"50",x"0d",x"0d",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"15",x"15",x"11",x"12",x"12",x"12",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"3a",x"3a",x"56",x"36",x"36",x"3a",x"3a",x"3a",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"36",x"36",x"3a",x"3a",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"33",x"33",x"33",x"33",x"33",x"13",x"12",x"12",x"33",x"33",x"33",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"56",x"79",x"98",x"75",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"76",x"d4",x"b4",x"d4",x"56",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"37",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"3b",x"3b",x"37",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"32",x"16",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"17",x"17",x"13",x"17",x"13",x"13",x"17",x"17",x"17",x"13",x"0e",x"12",x"17",x"13",x"12",x"13",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"37",x"12",x"12",x"12",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"16",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"37",x"3b",x"3b",x"37",x"17",x"17",x"17",x"37",x"37",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0a",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"12",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"99",x"b9",x"74",x"95",x"99",x"99",x"79",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"12",x"11",x"0d",x"0d",x"16",x"11",x"2c",x"2d",x"2d",x"2d",x"0d",x"0c",x"2d",x"2c",x"71",x"2c",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"12",x"12",x"12",x"11",x"11",x"16",x"16",x"12",x"12",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"56",x"36",x"36",x"3a",x"3a",x"3a",x"3a",x"3a",x"3a",x"3a",x"5a",x"3a",x"3a",x"36",x"36",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"13",x"33",x"33",x"33",x"37",x"33",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"75",x"99",x"98",x"55",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"b5",x"b4",x"b4",x"d4",x"56",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"37",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"3b",x"3b",x"3b",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"37",x"37",x"37",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"33",x"32",x"17",x"17",x"17",x"12",x"13",x"17",x"13",x"17",x"13",x"13",x"13",x"13",x"13",x"17",x"13",x"13",x"13",x"17",x"17",x"13",x"13",x"17",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"5b",x"37",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"16",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"37",x"3b",x"3b",x"37",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"56",x"99",x"95",x"51",x"55",x"79",x"79",x"79",x"79",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"51",x"11",x"0d",x"0d",x"16",x"2d",x"2c",x"2d",x"2d",x"2d",x"09",x"2d",x"2c",x"2d",x"51",x"2d",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"11",x"11",x"12",x"15",x"11",x"11",x"11",x"12",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"56",x"56",x"56",x"3a",x"3a",x"3a",x"3a",x"56",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"33",x"33",x"33",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0f",x"75",x"98",x"99",x"56",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"33",x"76",x"d8",x"b4",x"b4",x"d4",x"56",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"37",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"1b",x"1b",x"1b",x"1b",x"1b",x"3b",x"3b",x"1b",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"3b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"13",x"0e",x"12",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"13",x"13",x"17",x"17",x"13",x"12",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"12",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"17",x"17",x"3b",x"3b",x"37",x"17",x"17",x"17",x"37",x"37",x"17",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"55",x"75",x"51",x"51",x"51",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"55",x"55",x"55",x"55",x"55",x"31",x"0d",x"0d",x"12",x"2d",x"2c",x"2d",x"2d",x"0d",x"09",x"2d",x"2c",x"2d",x"2c",x"2d",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"12",x"11",x"11",x"11",x"11",x"11",x"15",x"16",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"5a",x"3a",x"3a",x"3a",x"3a",x"3a",x"3a",x"3a",x"36",x"36",x"36",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"79",x"98",x"95",x"56",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"13",x"13",x"13",x"76",x"f9",x"f8",x"b4",x"b4",x"f8",x"76",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"1b",x"1b",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"37",x"37",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"12",x"0e",x"12",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"13",x"0e",x"0e",x"12",x"12",x"17",x"17",x"13",x"0e",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"37",x"17",x"17",x"12",x"32",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"13",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"1b",x"37",x"3b",x"17",x"17",x"37",x"3b",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"56",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"55",x"75",x"51",x"4c",x"4c",x"51",x"75",x"75",x"75",x"51",x"51",x"51",x"55",x"55",x"55",x"75",x"31",x"0d",x"0d",x"11",x"2c",x"29",x"29",x"09",x"09",x"0d",x"2d",x"2c",x"2d",x"2c",x"0d",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"12",x"11",x"11",x"11",x"12",x"16",x"12",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"3a",x"3a",x"3a",x"5a",x"36",x"36",x"36",x"36",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"33",x"33",x"37",x"17",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"79",x"98",x"75",x"36",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"56",x"95",x"d8",x"f8",x"f8",x"b4",x"b4",x"f8",x"b9",x"37",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"37",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"37",x"37",x"37",x"37",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"37",x"37",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"17",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"12",x"13",x"12",x"0e",x"12",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"13",x"17",x"17",x"17",x"13",x"13",x"17",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"13",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"1b",x"17",x"17",x"17",x"17",x"1b",x"17",x"37",x"3b",x"1b",x"3b",x"3b",x"37",x"17",x"37",x"3b",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"95",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"55",x"75",x"71",x"51",x"50",x"2c",x"50",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"2d",x"0d",x"2d",x"29",x"29",x"2d",x"09",x"09",x"2d",x"2d",x"2c",x"2d",x"2c",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"12",x"12",x"15",x"11",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"33",x"13",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"32",x"79",x"98",x"75",x"32",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"32",x"95",x"f8",x"f8",x"f8",x"d8",x"94",x"b4",x"f8",x"f8",x"96",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"37",x"17",x"37",x"37",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"17",x"37",x"37",x"17",x"1b",x"1b",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"3b",x"37",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"13",x"12",x"12",x"12",x"0e",x"12",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"17",x"13",x"13",x"17",x"17",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"3b",x"37",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"17",x"17",x"1b",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"17",x"17",x"37",x"3b",x"17",x"17",x"17",x"37",x"17",x"17",x"37",x"37",x"1b",x"17",x"1b",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"16",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"b5",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"55",x"75",x"71",x"51",x"2d",x"31",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"0d",x"2d",x"29",x"29",x"0d",x"09",x"09",x"2d",x"2d",x"2c",x"2d",x"2d",x"09",x"09",x"09",x"0d",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"11",x"11",x"12",x"12",x"12",x"12",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"15",x"16",x"11",x"11",x"11",x"0d",x"0d",x"11",x"11",x"0d",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"3a",x"3a",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"33",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"56",x"95",x"98",x"75",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"95",x"f8",x"f8",x"f9",x"f9",x"d8",x"94",x"b4",x"f8",x"f8",x"d8",x"76",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"33",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"13",x"13",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"12",x"17",x"13",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"17",x"17",x"13",x"13",x"13",x"17",x"17",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"17",x"17",x"37",x"3b",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"3b",x"1b",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"12",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"75",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"75",x"36",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"75",x"95",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"51",x"71",x"51",x"51",x"51",x"2c",x"2d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"2d",x"29",x"29",x"2d",x"0d",x"09",x"29",x"2d",x"2d",x"2c",x"2c",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"11",x"11",x"12",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"12",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"12",x"12",x"11",x"11",x"12",x"16",x"36",x"36",x"36",x"36",x"36",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"55",x"99",x"98",x"55",x"13",x"13",x"13",x"12",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"d9",x"f8",x"f8",x"f9",x"f9",x"d8",x"94",x"b4",x"f9",x"f8",x"f8",x"b9",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"32",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"13",x"17",x"17",x"17",x"37",x"37",x"17",x"37",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"37",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"3b",x"37",x"3b",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"3b",x"17",x"17",x"37",x"3b",x"17",x"17",x"17",x"37",x"37",x"17",x"1b",x"1b",x"1b",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"11",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"95",x"d8",x"75",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"56",x"75",x"36",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"d5",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"31",x"51",x"51",x"51",x"51",x"2d",x"2d",x"2d",x"51",x"51",x"51",x"31",x"51",x"51",x"2d",x"29",x"2d",x"2d",x"08",x"09",x"29",x"2d",x"2d",x"2c",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"0d",x"0d",x"0e",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"16",x"36",x"36",x"36",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"75",x"79",x"98",x"56",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"f8",x"f8",x"f9",x"f9",x"f8",x"d8",x"94",x"d4",x"f9",x"fd",x"fc",x"d9",x"33",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"1b",x"17",x"17",x"1b",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"3b",x"37",x"37",x"3b",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"1b",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"1b",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"0d",x"11",x"12",x"16",x"15",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"16",x"16",x"16",x"16",x"16",x"d9",x"f8",x"d9",x"56",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"99",x"55",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"d1",x"72",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"31",x"51",x"51",x"51",x"51",x"2d",x"2d",x"2d",x"2d",x"4d",x"51",x"51",x"51",x"2d",x"29",x"29",x"09",x"09",x"29",x"29",x"2d",x"2d",x"2c",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"16",x"16",x"11",x"11",x"11",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"79",x"79",x"98",x"36",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"f8",x"f8",x"f9",x"f9",x"f8",x"d4",x"94",x"d4",x"f9",x"fd",x"fc",x"b9",x"37",x"17",x"17",x"17",x"13",x"17",x"13",x"0e",x"0e",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"13",x"13",x"12",x"12",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"12",x"17",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"17",x"37",x"37",x"3b",x"17",x"37",x"37",x"37",x"37",x"37",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"16",x"17",x"17",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"3b",x"1b",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"16",x"d4",x"f5",x"f9",x"9a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"75",x"95",x"36",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"d1",x"95",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"51",x"4d",x"51",x"51",x"2d",x"2c",x"2d",x"2d",x"4d",x"51",x"31",x"2d",x"29",x"29",x"09",x"29",x"29",x"29",x"2d",x"2d",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"0e",x"0e",x"0d",x"12",x"16",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"3a",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"99",x"78",x"98",x"36",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"d5",x"f8",x"f8",x"f8",x"f8",x"d4",x"94",x"b4",x"f9",x"fd",x"f8",x"b5",x"13",x"17",x"17",x"13",x"13",x"17",x"13",x"0e",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"13",x"13",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"13",x"13",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"37",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"16",x"16",x"f9",x"d5",x"f9",x"b9",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"55",x"95",x"55",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"d1",x"b5",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"2d",x"4d",x"4d",x"2d",x"2d",x"2c",x"2d",x"2d",x"2d",x"4d",x"2d",x"09",x"09",x"09",x"29",x"29",x"28",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"98",x"98",x"99",x"32",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"71",x"d4",x"f8",x"f8",x"d8",x"b4",x"b4",x"b4",x"d9",x"f8",x"f8",x"96",x"13",x"36",x"13",x"13",x"13",x"17",x"13",x"0e",x"12",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"13",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"3b",x"3b",x"3b",x"3b",x"3b",x"17",x"17",x"37",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"12",x"12",x"12",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"13",x"13",x"13",x"13",x"12",x"0e",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"37",x"17",x"37",x"37",x"17",x"17",x"37",x"37",x"37",x"37",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"16",x"16",x"f9",x"d5",x"f9",x"d9",x"76",x"16",x"3a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"1a",x"56",x"95",x"75",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"d1",x"d5",x"56",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"2d",x"4d",x"2d",x"2d",x"2c",x"2d",x"2d",x"2d",x"4d",x"2d",x"09",x"09",x"29",x"29",x"29",x"29",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3b",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"78",x"98",x"75",x"32",x"0f",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"72",x"d4",x"d8",x"b4",x"b4",x"b4",x"b4",x"d4",x"f8",x"b5",x"57",x"57",x"96",x"17",x"13",x"13",x"13",x"12",x"0e",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"17",x"3b",x"3b",x"1b",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"37",x"3b",x"3b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"37",x"37",x"17",x"17",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"16",x"76",x"f9",x"d5",x"d5",x"f9",x"b9",x"16",x"16",x"36",x"36",x"36",x"36",x"16",x"36",x"36",x"16",x"16",x"36",x"75",x"98",x"75",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"52",x"b5",x"d5",x"55",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"16",x"16",x"15",x"15",x"15",x"16",x"16",x"31",x"4d",x"4c",x"2d",x"2d",x"2c",x"2d",x"2d",x"2d",x"2d",x"09",x"09",x"29",x"29",x"29",x"29",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"3a",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"36",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"98",x"98",x"75",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"71",x"b5",x"b4",x"b4",x"b4",x"b4",x"d4",x"b5",x"56",x"56",x"d5",x"96",x"13",x"13",x"13",x"13",x"12",x"0e",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"13",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"17",x"37",x"37",x"3b",x"1b",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"13",x"13",x"12",x"12",x"12",x"13",x"17",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"32",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"37",x"3b",x"3b",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"16",x"16",x"d9",x"f9",x"b5",x"d5",x"f9",x"d9",x"56",x"1a",x"3a",x"3a",x"3a",x"3a",x"3a",x"3a",x"3a",x"1a",x"1a",x"1a",x"79",x"94",x"75",x"36",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"75",x"d1",x"d5",x"52",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"15",x"16",x"16",x"15",x"16",x"15",x"16",x"15",x"16",x"16",x"15",x"31",x"2d",x"4c",x"2c",x"2c",x"2d",x"2d",x"2d",x"2d",x"09",x"09",x"29",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"16",x"16",x"16",x"16",x"3a",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"36",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"98",x"98",x"75",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"95",x"b4",x"94",x"b4",x"b4",x"d4",x"76",x"37",x"96",x"f8",x"76",x"13",x"13",x"13",x"13",x"12",x"0e",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"0e",x"12",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"3b",x"3b",x"37",x"37",x"37",x"37",x"17",x"37",x"37",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"17",x"17",x"16",x"36",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"37",x"33",x"33",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"16",x"56",x"f9",x"f9",x"b5",x"d5",x"f9",x"f9",x"96",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"55",x"74",x"75",x"5a",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"95",x"d1",x"d5",x"52",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"15",x"15",x"16",x"16",x"15",x"15",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"31",x"2c",x"2c",x"2d",x"2d",x"2d",x"2d",x"2d",x"09",x"29",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"09",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"16",x"16",x"16",x"36",x"36",x"36",x"3a",x"36",x"36",x"36",x"36",x"1a",x"16",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"2e",x"2e",x"2e",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"98",x"98",x"55",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"91",x"d4",x"95",x"b4",x"d4",x"95",x"33",x"96",x"f8",x"f8",x"57",x"13",x"13",x"13",x"13",x"0e",x"0e",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"13",x"17",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"13",x"13",x"17",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"37",x"37",x"37",x"17",x"37",x"37",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"33",x"12",x"12",x"32",x"33",x"12",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"33",x"13",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"33",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"12",x"16",x"16",x"16",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"b5",x"f9",x"f9",x"b5",x"d5",x"f9",x"f9",x"b5",x"0e",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"52",x"75",x"74",x"99",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"b5",x"b1",x"d5",x"52",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"15",x"12",x"12",x"11",x"31",x"31",x"12",x"15",x"16",x"16",x"16",x"16",x"15",x"16",x"16",x"15",x"15",x"16",x"16",x"15",x"16",x"15",x"2c",x"2c",x"2c",x"2d",x"2d",x"2d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"0d",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"09",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"12",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"3a",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0a",x"0e",x"2e",x"51",x"51",x"75",x"75",x"75",x"75",x"75",x"55",x"51",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"55",x"78",x"78",x"55",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"95",x"d4",x"90",x"b4",x"d4",x"56",x"76",x"d9",x"f8",x"d9",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"37",x"17",x"17",x"37",x"17",x"37",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"13",x"13",x"32",x"13",x"17",x"17",x"37",x"33",x"17",x"17",x"13",x"17",x"17",x"17",x"13",x"32",x"33",x"13",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"33",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"13",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"12",x"13",x"17",x"17",x"17",x"16",x"16",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"f5",x"f9",x"f9",x"b5",x"d5",x"f9",x"f9",x"d5",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"51",x"94",x"79",x"36",x"16",x"16",x"12",x"12",x"12",x"12",x"32",x"f5",x"b1",x"d5",x"51",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"15",x"15",x"16",x"12",x"55",x"95",x"36",x"16",x"16",x"15",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"11",x"11",x"0d",x"09",x"2c",x"28",x"2d",x"4d",x"2d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"0e",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"11",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"2e",x"55",x"99",x"b8",x"b8",x"98",x"b8",x"b8",x"b8",x"b8",x"98",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"75",x"78",x"78",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"52",x"b5",x"b4",x"90",x"b4",x"b4",x"76",x"d9",x"fc",x"f8",x"b5",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"13",x"13",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"13",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"17",x"37",x"17",x"37",x"17",x"17",x"17",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"17",x"37",x"32",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"32",x"33",x"33",x"13",x"17",x"17",x"13",x"13",x"33",x"33",x"33",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"16",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"32",x"f9",x"f9",x"f9",x"b5",x"d5",x"f9",x"f9",x"d9",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"71",x"98",x"75",x"79",x"16",x"16",x"12",x"12",x"12",x"12",x"52",x"f5",x"b1",x"b5",x"56",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"12",x"15",x"15",x"15",x"16",x"75",x"b9",x"75",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"0d",x"0d",x"09",x"09",x"09",x"29",x"2c",x"4c",x"51",x"2d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"0e",x"0d",x"09",x"0d",x"0e",x"0d",x"0d",x"09",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"0d",x"09",x"09",x"09",x"09",x"0e",x"0a",x"2e",x"55",x"99",x"98",x"b8",x"98",x"98",x"75",x"75",x"99",x"98",x"b8",x"98",x"95",x"75",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"75",x"78",x"98",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"95",x"d4",x"b4",x"94",x"b4",x"b4",x"d9",x"d8",x"f8",x"f9",x"96",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"13",x"13",x"13",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"1b",x"17",x"37",x"37",x"17",x"37",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"37",x"17",x"17",x"17",x"32",x"33",x"33",x"13",x"13",x"33",x"32",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"16",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"51",x"f9",x"fd",x"f9",x"b5",x"d5",x"f9",x"fd",x"d5",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"98",x"51",x"99",x"16",x"16",x"16",x"16",x"12",x"12",x"96",x"f5",x"b1",x"b5",x"36",x"12",x"12",x"12",x"12",x"11",x"0d",x"11",x"11",x"0d",x"0d",x"11",x"16",x"15",x"15",x"16",x"75",x"b8",x"b9",x"75",x"16",x"16",x"16",x"16",x"11",x"11",x"0d",x"0d",x"09",x"09",x"09",x"05",x"05",x"05",x"09",x"09",x"70",x"70",x"2d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0a",x"2e",x"75",x"98",x"b8",x"99",x"75",x"51",x"31",x"32",x"32",x"32",x"51",x"75",x"99",x"b8",x"98",x"55",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"75",x"78",x"98",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"51",x"51",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"52",x"b5",x"d4",x"d4",x"b4",x"90",x"b4",x"b4",x"d8",x"d8",x"f8",x"d9",x"52",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"1b",x"37",x"37",x"37",x"37",x"37",x"17",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"13",x"12",x"13",x"12",x"12",x"13",x"17",x"13",x"12",x"17",x"13",x"13",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"31",x"f9",x"d9",x"f9",x"b5",x"d5",x"f9",x"f9",x"b5",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"95",x"54",x"98",x"36",x"16",x"16",x"16",x"16",x"36",x"d5",x"b1",x"d5",x"95",x"36",x"16",x"16",x"15",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"15",x"16",x"16",x"16",x"36",x"75",x"b9",x"b9",x"99",x"55",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"29",x"29",x"29",x"51",x"51",x"51",x"2c",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0e",x"75",x"98",x"98",x"75",x"51",x"0e",x"0a",x"0e",x"0e",x"0a",x"0a",x"0e",x"32",x"75",x"98",x"98",x"98",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"79",x"79",x"98",x"31",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"99",x"98",x"75",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"91",x"d8",x"f8",x"f8",x"d4",x"b4",x"b0",x"b5",x"d4",x"b4",x"d8",x"f8",x"d9",x"33",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"13",x"13",x"13",x"13",x"33",x"33",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"13",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"37",x"37",x"37",x"17",x"3b",x"1b",x"1b",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"12",x"0e",x"12",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"16",x"17",x"16",x"17",x"17",x"17",x"17",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"2e",x"b5",x"d5",x"d5",x"b5",x"b5",x"d5",x"d5",x"95",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"75",x"74",x"95",x"71",x"16",x"16",x"16",x"16",x"56",x"f5",x"b1",x"f5",x"96",x"16",x"16",x"16",x"15",x"15",x"15",x"15",x"15",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"75",x"b9",x"95",x"b8",x"b9",x"51",x"09",x"05",x"09",x"29",x"29",x"2d",x"2d",x"4d",x"4d",x"51",x"51",x"71",x"95",x"95",x"0d",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"75",x"98",x"98",x"75",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"75",x"b8",x"98",x"95",x"2e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"78",x"74",x"98",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"95",x"98",x"51",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"d5",x"d8",x"f8",x"f8",x"f8",x"d4",x"94",x"b4",x"b4",x"d4",x"d8",x"fc",x"f8",x"b5",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"13",x"33",x"52",x"71",x"91",x"b5",x"b1",x"72",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"13",x"13",x"12",x"0e",x"12",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"16",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"16",x"16",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"71",x"d5",x"d5",x"95",x"b5",x"d5",x"b5",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"75",x"98",x"55",x"95",x"0d",x"0e",x"12",x"36",x"96",x"f5",x"b1",x"f5",x"56",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"0d",x"09",x"09",x"51",x"b8",x"b8",x"b8",x"b8",x"b8",x"94",x"b5",x"b8",x"b8",x"b8",x"b8",x"b8",x"94",x"74",x"94",x"b8",x"98",x"51",x"2d",x"09",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"11",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"2d",x"99",x"98",x"75",x"2e",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"31",x"95",x"98",x"98",x"51",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"98",x"74",x"98",x"32",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"75",x"99",x"75",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"91",x"f8",x"f8",x"d8",x"d8",x"f8",x"b4",x"94",x"b4",x"d4",x"d8",x"d8",x"f8",x"f8",x"96",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"2e",x"72",x"92",x"b1",x"d1",x"d5",x"d5",x"d1",x"ad",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"12",x"0e",x"0e",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"13",x"13",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"16",x"16",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"95",x"b5",x"b5",x"b5",x"b5",x"91",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"51",x"98",x"51",x"b8",x"2d",x"0e",x"0e",x"32",x"d5",x"d1",x"d5",x"d5",x"36",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"2d",x"71",x"b8",x"94",x"94",x"94",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"bc",x"bc",x"b8",x"98",x"95",x"75",x"51",x"2d",x"09",x"09",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"2d",x"75",x"98",x"75",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"98",x"98",x"99",x"51",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"78",x"75",x"78",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"75",x"98",x"51",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"d5",x"f8",x"d8",x"d8",x"d8",x"f8",x"b4",x"90",x"b4",x"d8",x"d8",x"d8",x"f8",x"f9",x"76",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"6e",x"cd",x"f1",x"d5",x"d5",x"d5",x"b1",x"b1",x"cd",x"4e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"16",x"16",x"16",x"17",x"16",x"17",x"17",x"17",x"17",x"16",x"17",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"0d",x"09",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"52",x"b5",x"b5",x"b5",x"95",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"98",x"30",x"98",x"51",x"0e",x"0a",x"6d",x"d5",x"91",x"f9",x"91",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"05",x"09",x"09",x"4d",x"95",x"b8",x"98",x"74",x"75",x"70",x"95",x"94",x"74",x"75",x"74",x"94",x"98",x"98",x"b8",x"95",x"71",x"2d",x"09",x"09",x"09",x"09",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"0d",x"0e",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"11",x"11",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"1a",x"1a",x"1a",x"1a",x"1a",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"51",x"98",x"98",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"12",x"75",x"98",x"98",x"75",x"32",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"36",x"78",x"74",x"78",x"36",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"75",x"99",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"52",x"f8",x"d8",x"f8",x"d8",x"d8",x"d8",x"b4",x"90",x"b4",x"d8",x"d8",x"d8",x"f8",x"d5",x"72",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"32",x"52",x"32",x"52",x"b1",x"ad",x"8d",x"ad",x"52",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"16",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"16",x"17",x"17",x"17",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"b5",x"b5",x"b5",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"31",x"99",x"55",x"98",x"75",x"0e",x"2e",x"91",x"d5",x"b1",x"f9",x"4d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"4d",x"71",x"74",x"75",x"94",x"94",x"98",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"94",x"71",x"4d",x"2d",x"29",x"09",x"09",x"09",x"09",x"0d",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"2d",x"75",x"98",x"51",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"55",x"99",x"98",x"99",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"55",x"74",x"74",x"74",x"36",x"16",x"1a",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"0e",x"51",x"b8",x"75",x"0e",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"52",x"f8",x"f8",x"f9",x"d8",x"d8",x"d8",x"b4",x"90",x"b4",x"f8",x"d8",x"d8",x"f8",x"d4",x"72",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"92",x"ad",x"89",x"8d",x"32",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"12",x"12",x"13",x"13",x"13",x"12",x"0e",x"0e",x"12",x"13",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"13",x"12",x"17",x"17",x"17",x"13",x"32",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"b5",x"b5",x"b5",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"99",x"75",x"75",x"99",x"2d",x"52",x"b5",x"b1",x"d5",x"d5",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"71",x"98",x"98",x"98",x"98",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"95",x"51",x"09",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"0d",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"51",x"b8",x"95",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"79",x"98",x"98",x"79",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"55",x"74",x"75",x"74",x"35",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"98",x"98",x"32",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"b5",x"f8",x"d9",x"d9",x"d8",x"d8",x"b4",x"90",x"d4",x"f8",x"d8",x"d8",x"d8",x"d4",x"71",x"0e",x"13",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"13",x"13",x"13",x"13",x"52",x"8d",x"89",x"6d",x"33",x"13",x"12",x"12",x"13",x"13",x"12",x"13",x"12",x"13",x"13",x"0e",x"12",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"13",x"32",x"16",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"13",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"17",x"17",x"17",x"17",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"0e",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"d5",x"d5",x"b5",x"b5",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"2e",x"75",x"99",x"55",x"b8",x"51",x"92",x"d5",x"b1",x"f9",x"91",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"95",x"75",x"94",x"b8",x"dc",x"dc",x"b8",x"b8",x"94",x"94",x"99",x"99",x"75",x"75",x"75",x"75",x"51",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"08",x"08",x"09",x"09",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"75",x"98",x"51",x"05",x"09",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"15",x"12",x"55",x"98",x"b8",x"99",x"35",x"16",x"12",x"11",x"12",x"12",x"11",x"55",x"74",x"75",x"74",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"79",x"b8",x"59",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"71",x"d8",x"d8",x"d8",x"d8",x"b4",x"94",x"90",x"b4",x"f9",x"d8",x"d9",x"d8",x"d8",x"91",x"0e",x"0e",x"12",x"13",x"13",x"0e",x"0e",x"0e",x"13",x"13",x"13",x"13",x"32",x"8d",x"88",x"6d",x"32",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"16",x"12",x"12",x"12",x"17",x"13",x"12",x"12",x"12",x"12",x"13",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"b5",x"f9",x"b4",x"90",x"d5",x"95",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"75",x"b8",x"31",x"98",x"95",x"b1",x"d1",x"d5",x"f5",x"2d",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"51",x"94",x"b8",x"d8",x"b9",x"95",x"4d",x"4d",x"75",x"50",x"4c",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"99",x"75",x"09",x"09",x"0d",x"15",x"15",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"11",x"12",x"35",x"79",x"b8",x"98",x"75",x"12",x"12",x"11",x"11",x"12",x"11",x"55",x"75",x"75",x"75",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"98",x"98",x"36",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"b4",x"d4",x"b4",x"b4",x"b4",x"90",x"90",x"b4",x"d9",x"d9",x"d9",x"d8",x"f8",x"95",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"13",x"13",x"12",x"13",x"52",x"6d",x"69",x"6d",x"4e",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"13",x"17",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"16",x"16",x"15",x"11",x"11",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"51",x"b5",x"f9",x"f8",x"b0",x"90",x"f4",x"d5",x"52",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"b8",x"31",x"98",x"d9",x"b1",x"b1",x"f9",x"b5",x"09",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"51",x"98",x"98",x"b8",x"94",x"71",x"2d",x"09",x"09",x"51",x"51",x"2c",x"50",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"09",x"05",x"09",x"09",x"0d",x"09",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"31",x"2d",x"2d",x"11",x"11",x"11",x"0d"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"75",x"b8",x"51",x"05",x"0d",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"12",x"12",x"16",x"59",x"98",x"98",x"99",x"12",x"12",x"11",x"11",x"12",x"12",x"55",x"75",x"75",x"75",x"11",x"12",x"16",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"75",x"b8",x"75",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"b4",x"b4",x"b4",x"94",x"90",x"90",x"b4",x"b4",x"d4",x"d8",x"d8",x"d8",x"b5",x"4e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"13",x"13",x"12",x"13",x"4e",x"8d",x"69",x"69",x"6d",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"13",x"17",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"17",x"17",x"17",x"17",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0a",x"71",x"d9",x"f9",x"f9",x"f8",x"90",x"90",x"d4",x"f8",x"b5",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2d",x"b8",x"55",x"95",x"b5",x"b1",x"d5",x"d5",x"4e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"94",x"dc",x"b8",x"51",x"09",x"05",x"09",x"09",x"09",x"2d",x"75",x"50",x"2c",x"50",x"75",x"75",x"75",x"75",x"54",x"75",x"74",x"2d",x"05",x"09",x"09",x"0d",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"05",x"09",x"2d",x"2c",x"50",x"50",x"30",x"50",x"74",x"74",x"75",x"75",x"75",x"51",x"51"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"95",x"95",x"2d",x"0d",x"15",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"16",x"16",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"16",x"59",x"99",x"98",x"99",x"51",x"12",x"11",x"11",x"12",x"12",x"55",x"75",x"75",x"75",x"11",x"12",x"12",x"11",x"12",x"12",x"16",x"16",x"16",x"12",x"35",x"99",x"b8",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"95",x"b4",x"94",x"90",x"90",x"90",x"94",x"b4",x"b4",x"b4",x"d8",x"d4",x"b4",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"6d",x"6d",x"69",x"69",x"8d",x"6d",x"72",x"52",x"32",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"13",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"13",x"13",x"17",x"17",x"17",x"17",x"12",x"12",x"17",x"12",x"12",x"12",x"13",x"17",x"17",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"b5",x"fd",x"f9",x"f8",x"f8",x"90",x"90",x"d4",x"f8",x"d9",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"b8",x"74",x"95",x"b1",x"d5",x"d5",x"b5",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"2d",x"95",x"b8",x"95",x"2d",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"50",x"50",x"2c",x"4c",x"51",x"55",x"75",x"75",x"55",x"55",x"75",x"51",x"09",x"05",x"09",x"09",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"2d",x"2d",x"2c",x"50",x"51",x"30",x"50",x"50",x"74",x"74",x"70",x"51",x"71",x"75"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"99",x"75",x"0d",x"12",x"16",x"16",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"16",x"35",x"75",x"98",x"99",x"75",x"12",x"12",x"11",x"12",x"11",x"55",x"75",x"75",x"75",x"11",x"12",x"11",x"11",x"12",x"12",x"16",x"12",x"12",x"12",x"55",x"b8",x"95",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"71",x"90",x"90",x"90",x"90",x"91",x"90",x"b4",x"b4",x"b4",x"b4",x"b4",x"90",x"90",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"8d",x"69",x"69",x"8d",x"ac",x"8d",x"8d",x"72",x"52",x"32",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"13",x"0e",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"12",x"12",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"2d",x"d5",x"fd",x"d9",x"f8",x"f8",x"90",x"90",x"d8",x"f8",x"f9",x"b5",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"99",x"94",x"b5",x"b1",x"d5",x"d5",x"71",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"75",x"b8",x"95",x"2d",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"2c",x"50",x"4c",x"2c",x"50",x"51",x"50",x"55",x"55",x"51",x"51",x"75",x"2d",x"09",x"09",x"09",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"2c",x"2c",x"2c",x"2c",x"2c",x"2d",x"2c",x"2c",x"2c",x"51",x"50",x"50",x"50",x"71",x"74"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"51",x"99",x"55",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"12",x"12",x"11",x"12",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"12",x"16",x"12",x"55",x"98",x"99",x"98",x"12",x"12",x"11",x"11",x"11",x"75",x"75",x"75",x"75",x"11",x"12",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"35",x"95",x"b8",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"52",x"90",x"90",x"90",x"90",x"91",x"90",x"91",x"b4",x"b4",x"b4",x"90",x"90",x"90",x"4d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4d",x"8d",x"8d",x"8d",x"69",x"69",x"69",x"69",x"69",x"b1",x"d5",x"b1",x"52",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"13",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"13",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"4e",x"d5",x"f8",x"d8",x"f8",x"f8",x"90",x"b0",x"d8",x"f8",x"f8",x"b5",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"75",x"98",x"d5",x"b1",x"d5",x"b5",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"05",x"51",x"b8",x"94",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"50",x"51",x"2c",x"2c",x"51",x"51",x"50",x"54",x"54",x"51",x"51",x"51",x"09",x"09",x"09",x"08",x"08",x"09",x"09",x"09",x"09",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"08",x"08",x"2c",x"30",x"54",x"74",x"74"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"75",x"99",x"35",x"16",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"12",x"12",x"12",x"35",x"98",x"98",x"98",x"31",x"11",x"12",x"12",x"11",x"75",x"75",x"75",x"75",x"11",x"12",x"11",x"11",x"12",x"12",x"12",x"11",x"12",x"55",x"b8",x"99",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"91",x"90",x"90",x"90",x"91",x"90",x"95",x"b4",x"b4",x"b4",x"94",x"90",x"90",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"6d",x"ad",x"ad",x"ad",x"ad",x"8d",x"8d",x"89",x"8d",x"b1",x"d5",x"d5",x"96",x"13",x"13",x"13",x"12",x"13",x"13",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"16",x"12",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"16",x"12",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"b5",x"f8",x"f8",x"f8",x"d8",x"90",x"b0",x"d8",x"fc",x"f8",x"95",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"75",x"b9",x"b1",x"d5",x"f5",x"91",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"4d",x"b8",x"99",x"4d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"50",x"50",x"2c",x"4c",x"50",x"50",x"50",x"51",x"51",x"51",x"51",x"2d",x"05",x"09",x"08",x"09",x"09",x"09",x"09",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"08",x"08",x"08",x"2c",x"4c",x"51",x"75",x"74",x"74",x"50"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"98",x"99",x"35",x"11",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"12",x"31",x"95",x"98",x"98",x"75",x"12",x"12",x"12",x"11",x"75",x"75",x"74",x"55",x"11",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"75",x"b8",x"75",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"91",x"90",x"90",x"90",x"91",x"90",x"b4",x"b4",x"b4",x"b4",x"b4",x"90",x"90",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4d",x"ad",x"ad",x"ad",x"cd",x"ad",x"ad",x"ad",x"b1",x"91",x"b1",x"d5",x"d1",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"16",x"12",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"3a",x"3a",x"3a",x"3a",x"3a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"71",x"d4",x"f4",x"d4",x"b4",x"90",x"90",x"d4",x"f8",x"d4",x"71",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"d9",x"b1",x"d5",x"f9",x"75",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"95",x"b8",x"51",x"09",x"09",x"09",x"09",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"50",x"51",x"4c",x"2c",x"50",x"51",x"4c",x"51",x"51",x"51",x"51",x"2d",x"05",x"08",x"08",x"09",x"09",x"09",x"2c",x"2c",x"2c",x"28",x"28",x"28",x"28",x"2c",x"08",x"08",x"2c",x"50",x"74",x"95",x"75",x"75",x"51",x"2d"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"31",x"98",x"75",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"12",x"12",x"75",x"98",x"98",x"99",x"12",x"12",x"12",x"11",x"75",x"75",x"75",x"55",x"11",x"12",x"12",x"11",x"11",x"12",x"11",x"12",x"31",x"95",x"98",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"91",x"90",x"90",x"90",x"90",x"91",x"90",x"b4",x"d8",x"d4",x"b4",x"b4",x"b0",x"90",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"8d",x"d1",x"d1",x"d1",x"b1",x"b1",x"b5",x"d5",x"b1",x"b1",x"d1",x"cd",x"33",x"12",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"17",x"12",x"12",x"12",x"17",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"16",x"16",x"16",x"16",x"11",x"11",x"12",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"09",x"09",x"4d",x"b4",x"d4",x"90",x"90",x"b0",x"b0",x"d4",x"b1",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"31",x"d9",x"b1",x"d5",x"d9",x"75",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"2d",x"d8",x"74",x"0d",x"09",x"09",x"09",x"2d",x"95",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"50",x"50",x"2c",x"2c",x"51",x"50",x"4c",x"51",x"51",x"50",x"2d",x"05",x"08",x"08",x"09",x"09",x"2c",x"2c",x"2c",x"28",x"2c",x"2c",x"08",x"08",x"08",x"2c",x"50",x"75",x"74",x"74",x"75",x"75",x"51",x"0d",x"0d"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"11",x"35",x"b8",x"55",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"55",x"98",x"98",x"98",x"31",x"12",x"12",x"11",x"75",x"75",x"75",x"55",x"11",x"12",x"12",x"11",x"12",x"11",x"11",x"12",x"55",x"b8",x"98",x"31",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"71",x"b4",x"b4",x"90",x"90",x"90",x"91",x"94",x"d4",x"f8",x"f8",x"d4",x"b4",x"b4",x"90",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"b1",x"d1",x"d1",x"d5",x"d5",x"d5",x"91",x"8d",x"cd",x"ad",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"17",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"13",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"16",x"16",x"16",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"6d",x"b4",x"90",x"90",x"b0",x"b0",x"90",x"4d",x"09",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"b5",x"d5",x"d5",x"b9",x"75",x"2d",x"0e",x"0e",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"95",x"b8",x"2d",x"09",x"09",x"09",x"09",x"51",x"b9",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2c",x"50",x"2c",x"2c",x"2c",x"51",x"4c",x"50",x"50",x"50",x"31",x"09",x"08",x"08",x"09",x"28",x"2c",x"2c",x"28",x"28",x"28",x"08",x"08",x"0c",x"2c",x"2c",x"50",x"75",x"74",x"74",x"51",x"31",x"0d",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0d",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"11",x"11",x"12",x"12",x"55",x"99",x"31",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"12",x"11",x"12",x"31",x"98",x"98",x"98",x"55",x"11",x"12",x"11",x"75",x"75",x"75",x"55",x"11",x"12",x"11",x"12",x"12",x"11",x"12",x"12",x"75",x"b8",x"75",x"12",x"11",x"11",x"16",x"16",x"16",x"16",x"16",x"15",x"16",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"91",x"d8",x"d8",x"b4",x"90",x"90",x"90",x"94",x"b4",x"d4",x"f8",x"f8",x"d4",x"b4",x"b4",x"90",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4e",x"91",x"d1",x"d1",x"d1",x"b1",x"8d",x"69",x"ad",x"8d",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"17",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"1a",x"1a",x"1a",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"0e",x"0e",x"0e",x"12",x"0d",x"0d",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"29",x"b4",x"90",x"90",x"b0",x"b0",x"4d",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"91",x"f5",x"95",x"99",x"99",x"51",x"0e",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"2d",x"dc",x"74",x"09",x"09",x"09",x"09",x"09",x"95",x"dd",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"4c",x"50",x"2c",x"2c",x"4d",x"2c",x"2c",x"50",x"51",x"31",x"08",x"08",x"08",x"28",x"28",x"28",x"28",x"28",x"08",x"08",x"08",x"08",x"2c",x"2c",x"2c",x"50",x"70",x"70",x"51",x"2d",x"0d",x"09",x"0d",x"0d"),
(x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"55",x"99",x"31",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"12",x"11",x"11",x"12",x"11",x"99",x"98",x"98",x"75",x"11",x"12",x"31",x"75",x"75",x"75",x"55",x"11",x"12",x"12",x"11",x"12",x"11",x"12",x"31",x"95",x"b8",x"75",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"95",x"d8",x"d8",x"d8",x"d8",x"b4",x"90",x"90",x"94",x"b4",x"b4",x"d8",x"d8",x"f8",x"d4",x"d4",x"b4",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"ad",x"ad",x"ad",x"6d",x"69",x"8d",x"4e",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"12",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"0d",x"12",x"0e",x"0e",x"0d",x"12",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"09",x"09",x"29",x"b0",x"90",x"90",x"b4",x"6d",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"91",x"f5",x"75",x"74",x"b9",x"75",x"0a",x"0e",x"0e",x"0d",x"09",x"09",x"0d",x"95",x"98",x"51",x"09",x"09",x"09",x"09",x"0d",x"b9",x"bd",x"51",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"2c",x"4c",x"31",x"2c",x"2c",x"2c",x"2c",x"2c",x"50",x"50",x"08",x"08",x"08",x"28",x"28",x"29",x"28",x"08",x"08",x"08",x"08",x"2c",x"2c",x"2c",x"2c",x"4c",x"4c",x"2c",x"0d",x"09",x"09",x"0d",x"0d",x"0d"),
(x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"75",x"75",x"31",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"12",x"11",x"75",x"98",x"98",x"99",x"31",x"12",x"31",x"74",x"75",x"75",x"55",x"11",x"12",x"12",x"12",x"12",x"16",x"16",x"55",x"99",x"98",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"52",x"95",x"d4",x"f8",x"d8",x"d8",x"d8",x"b4",x"90",x"90",x"b4",x"b4",x"d8",x"d8",x"d8",x"f8",x"f8",x"d4",x"71",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"8d",x"8d",x"69",x"69",x"6d",x"6d",x"32",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"12",x"12",x"13",x"12",x"13",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"12",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"12",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"4d",x"b4",x"90",x"b0",x"b4",x"4d",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"b1",x"f5",x"51",x"54",x"b9",x"95",x"0a",x"0e",x"0e",x"0d",x"09",x"09",x"2d",x"98",x"54",x"2d",x"09",x"09",x"09",x"09",x"4d",x"bc",x"b9",x"95",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"4c",x"2c",x"2c",x"2c",x"2c",x"2d",x"2c",x"4c",x"30",x"08",x"08",x"28",x"28",x"28",x"28",x"08",x"08",x"08",x"08",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d"),
(x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"95",x"75",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"55",x"98",x"99",x"99",x"31",x"12",x"31",x"74",x"75",x"75",x"55",x"11",x"12",x"12",x"12",x"12",x"16",x"16",x"75",x"98",x"79",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"91",x"b5",x"d8",x"d8",x"d8",x"d8",x"d8",x"d8",x"b4",x"70",x"90",x"b4",x"d8",x"d8",x"d8",x"d8",x"f8",x"f8",x"b5",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"6d",x"8d",x"69",x"69",x"6d",x"6d",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"12",x"12",x"13",x"12",x"12",x"13",x"12",x"12",x"12",x"12",x"17",x"13",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"16",x"1a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"0d",x"12",x"11",x"0d",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"29",x"6c",x"b4",x"90",x"b0",x"b0",x"2d",x"09",x"09",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"d5",x"d5",x"55",x"54",x"98",x"95",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"51",x"98",x"51",x"09",x"09",x"09",x"09",x"09",x"71",x"b8",x"95",x"99",x"2d",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"4c",x"2c",x"2c",x"2c",x"2c",x"2d",x"2d",x"2c",x"2c",x"08",x"08",x"28",x"28",x"28",x"08",x"08",x"08",x"28",x"28",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11"),
(x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"0d",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"95",x"55",x"11",x"12",x"11",x"11",x"12",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"55",x"55",x"31",x"0e",x"12",x"11",x"11",x"11",x"11",x"11",x"31",x"98",x"99",x"b8",x"55",x"12",x"31",x"75",x"75",x"75",x"55",x"11",x"12",x"11",x"11",x"11",x"12",x"16",x"79",x"b8",x"75",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"52",x"d8",x"d9",x"d8",x"d8",x"d8",x"d8",x"d8",x"d8",x"d8",x"94",x"70",x"90",x"b8",x"d8",x"d8",x"d8",x"d8",x"b5",x"52",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"6d",x"6d",x"69",x"69",x"6d",x"4d",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"12",x"12",x"13",x"13",x"12",x"13",x"12",x"12",x"12",x"12",x"17",x"13",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"12",x"0e",x"0e",x"11",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"05",x"09",x"4d",x"b4",x"d4",x"b0",x"70",x"b0",x"90",x"29",x"09",x"09",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"d5",x"d9",x"75",x"55",x"98",x"99",x"2d",x"0e",x"0e",x"0d",x"09",x"2d",x"71",x"50",x"50",x"09",x"09",x"09",x"05",x"2d",x"95",x"99",x"95",x"98",x"51",x"09",x"09",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"2d",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"0c",x"08",x"28",x"08",x"08",x"08",x"08",x"28",x"28",x"28",x"2c",x"2c",x"2c",x"2c",x"2c",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11"),
(x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"98",x"55",x"11",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"55",x"75",x"75",x"55",x"11",x"12",x"11",x"11",x"11",x"11",x"31",x"98",x"98",x"98",x"75",x"12",x"15",x"75",x"75",x"75",x"55",x"16",x"12",x"12",x"12",x"11",x"12",x"16",x"99",x"b8",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"0d",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"91",x"f8",x"fc",x"d8",x"d8",x"d8",x"d8",x"d8",x"d8",x"d8",x"90",x"70",x"94",x"d8",x"d8",x"d8",x"d8",x"d8",x"b5",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"6d",x"69",x"49",x"69",x"6d",x"32",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"12",x"12",x"13",x"17",x"13",x"12",x"13",x"12",x"12",x"12",x"12",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"1a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"12",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"29",x"6d",x"b4",x"f8",x"f4",x"90",x"70",x"b0",x"b4",x"29",x"05",x"09",x"0e",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"2d",x"f9",x"b5",x"75",x"55",x"74",x"b9",x"51",x"0a",x"0e",x"0d",x"09",x"2d",x"74",x"31",x"51",x"09",x"09",x"09",x"05",x"2d",x"b9",x"99",x"95",x"98",x"75",x"2d",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"11",x"11",x"0d",x"2d",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"0c",x"08",x"08",x"08",x"08",x"08",x"28",x"28",x"28",x"2c",x"2c",x"2c",x"2c",x"2d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d"),
(x"12",x"12",x"12",x"12",x"0d",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"98",x"55",x"11",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"55",x"95",x"b8",x"55",x"11",x"11",x"11",x"11",x"12",x"12",x"99",x"98",x"98",x"79",x"36",x"15",x"74",x"75",x"74",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"55",x"99",x"98",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"0d",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"d4",x"f8",x"d8",x"d8",x"d8",x"d9",x"d9",x"d9",x"d9",x"d8",x"90",x"70",x"b4",x"d8",x"d8",x"d8",x"d8",x"d8",x"d8",x"52",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4d",x"6d",x"6d",x"6d",x"69",x"69",x"8d",x"6d",x"2e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"13",x"17",x"13",x"12",x"13",x"12",x"12",x"12",x"12",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"12",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"b0",x"f8",x"f8",x"d8",x"d4",x"b0",x"90",x"b0",x"d4",x"4d",x"05",x"09",x"0e",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"4d",x"d5",x"b5",x"95",x"55",x"74",x"b8",x"75",x"09",x"0e",x"09",x"09",x"2d",x"50",x"51",x"31",x"09",x"09",x"09",x"09",x"51",x"bc",x"99",x"74",x"98",x"99",x"31",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"2d",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"08",x"08",x"08",x"08",x"08",x"28",x"28",x"08",x"28",x"2c",x"2c",x"2c",x"2c",x"0d",x"12",x"11",x"0d",x"11",x"0d",x"11",x"11",x"11",x"11",x"0d"),
(x"12",x"12",x"12",x"12",x"0d",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"95",x"31",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"31",x"75",x"98",x"55",x"11",x"11",x"11",x"12",x"12",x"75",x"98",x"98",x"99",x"35",x"11",x"74",x"55",x"74",x"55",x"16",x"16",x"15",x"16",x"16",x"16",x"75",x"98",x"98",x"55",x"16",x"16",x"16",x"16",x"12",x"0d",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"d8",x"f8",x"d9",x"d8",x"d8",x"d8",x"d8",x"d8",x"d8",x"b4",x"70",x"70",x"b4",x"d8",x"d8",x"d8",x"d9",x"d8",x"d8",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4e",x"8d",x"8d",x"8d",x"8d",x"69",x"49",x"6d",x"ad",x"8d",x"4e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"13",x"17",x"13",x"12",x"13",x"12",x"12",x"12",x"12",x"17",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"0d",x"0e",x"0e",x"0d",x"0d",x"09",x"70",x"d4",x"f8",x"d4",x"d4",x"d4",x"90",x"70",x"b4",x"f8",x"91",x"29",x"09",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"72",x"d5",x"95",x"99",x"55",x"54",x"b8",x"95",x"09",x"0d",x"09",x"09",x"2d",x"50",x"75",x"2d",x"09",x"09",x"09",x"0d",x"75",x"b8",x"95",x"71",x"99",x"98",x"55",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"2c",x"2c",x"28",x"2c",x"2d",x"2c",x"08",x"08",x"08",x"08",x"28",x"28",x"28",x"28",x"28",x"2c",x"2c",x"2d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"11",x"11",x"12",x"12",x"12",x"12"),
(x"12",x"12",x"12",x"12",x"0d",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"2d",x"51",x"2d",x"32",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"31",x"99",x"99",x"31",x"12",x"11",x"11",x"12",x"55",x"98",x"98",x"98",x"55",x"11",x"74",x"55",x"75",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"75",x"98",x"79",x"35",x"16",x"16",x"16",x"12",x"0d",x"09",x"09",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"d8",x"f8",x"f9",x"d8",x"b4",x"d8",x"d8",x"d8",x"d8",x"b4",x"70",x"70",x"b4",x"d8",x"d8",x"d8",x"d9",x"d8",x"d8",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"6d",x"ad",x"ad",x"ad",x"ad",x"8d",x"69",x"69",x"8d",x"ad",x"8e",x"32",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"13",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"b4",x"f8",x"d4",x"d4",x"d4",x"d4",x"90",x"70",x"d4",x"f8",x"d4",x"6d",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"92",x"b1",x"95",x"b9",x"75",x"51",x"b8",x"99",x"0d",x"0d",x"09",x"2d",x"2d",x"50",x"75",x"0d",x"09",x"0d",x"0d",x"31",x"99",x"b9",x"99",x"51",x"99",x"99",x"75",x"31",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"2c",x"2c",x"28",x"2c",x"2d",x"2c",x"08",x"08",x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"2d",x"2d",x"0d",x"0d",x"12",x"11",x"12",x"11",x"0d",x"11",x"16",x"16",x"16",x"16",x"16"),
(x"12",x"12",x"12",x"12",x"0d",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"2e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"2e",x"4d",x"4e",x"4e",x"4d",x"31",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"31",x"98",x"75",x"31",x"11",x"11",x"11",x"51",x"98",x"98",x"98",x"55",x"31",x"75",x"55",x"75",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"79",x"98",x"79",x"36",x"16",x"16",x"0d",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"d4",x"f8",x"f9",x"d8",x"b4",x"b4",x"d8",x"d8",x"b8",x"90",x"6c",x"90",x"b4",x"d8",x"d8",x"d8",x"d9",x"b8",x"d8",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"8d",x"ad",x"ad",x"ad",x"ad",x"ad",x"8d",x"69",x"49",x"ad",x"ad",x"91",x"32",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"13",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"12",x"0e",x"12",x"0d",x"0d",x"09",x"09",x"d5",x"d8",x"d8",x"d8",x"d8",x"d4",x"70",x"90",x"d4",x"d4",x"f8",x"b4",x"51",x"0e",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"91",x"b1",x"95",x"b9",x"75",x"51",x"98",x"b8",x"2d",x"0d",x"0d",x"31",x"50",x"50",x"75",x"0d",x"0d",x"0d",x"0d",x"51",x"b9",x"b9",x"99",x"51",x"99",x"99",x"78",x"51",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"11",x"16",x"12",x"2d",x"2c",x"2c",x"2c",x"2c",x"28",x"08",x"28",x"28",x"28",x"28",x"28",x"28",x"09",x"0d",x"0d",x"12",x"12",x"0d",x"11",x"16",x"16",x"11",x"11",x"11",x"15",x"15",x"11",x"16",x"16"),
(x"0e",x"12",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"2e",x"4e",x"4e",x"4e",x"4e",x"4d",x"4e",x"2e",x"4d",x"4d",x"49",x"2d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"75",x"98",x"55",x"12",x"11",x"11",x"31",x"99",x"99",x"98",x"75",x"35",x"74",x"75",x"75",x"55",x"15",x"16",x"16",x"16",x"16",x"35",x"78",x"98",x"55",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"b4",x"d8",x"d8",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"70",x"6c",x"90",x"b4",x"d8",x"d8",x"d8",x"d8",x"d8",x"f8",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"ad",x"ad",x"8d",x"8d",x"8d",x"8d",x"ad",x"8d",x"49",x"69",x"ad",x"d1",x"92",x"32",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"13",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"12",x"0e",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"13",x"13",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"0e",x"12",x"0e",x"12",x"0d",x"0d",x"09",x"09",x"b4",x"d8",x"d8",x"d8",x"d8",x"b4",x"6c",x"90",x"d8",x"d4",x"d4",x"d8",x"95",x"0e",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0d",x"0e",x"0e",x"0d",x"0e",x"0d",x"0d",x"0d",x"95",x"91",x"91",x"99",x"74",x"55",x"99",x"b8",x"51",x"0e",x"0e",x"31",x"50",x"50",x"75",x"0d",x"0d",x"0d",x"0d",x"55",x"b9",x"99",x"95",x"50",x"99",x"99",x"98",x"55",x"11",x"11",x"11",x"12",x"12",x"16",x"0d",x"0d",x"16",x"12",x"0d",x"2d",x"2c",x"2c",x"2c",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"16",x"12",x"12",x"11",x"12",x"16",x"16",x"16",x"16",x"16"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"2e",x"2e",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"4e",x"2e",x"2e",x"2d",x"2d",x"4d",x"4d",x"4e",x"4e",x"4d",x"4d",x"49",x"29",x"2d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"98",x"75",x"11",x"12",x"12",x"11",x"99",x"98",x"98",x"79",x"55",x"54",x"75",x"75",x"55",x"15",x"16",x"16",x"16",x"16",x"55",x"78",x"98",x"51",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2d",x"b0",x"d4",x"b4",x"b4",x"b9",x"b4",x"94",x"94",x"91",x"70",x"6c",x"70",x"b4",x"d8",x"b8",x"b8",x"d4",x"d8",x"f8",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"8d",x"b1",x"b1",x"ad",x"ad",x"8d",x"ad",x"ad",x"6d",x"49",x"8d",x"d1",x"d1",x"72",x"13",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"12",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"0d",x"0d",x"0d",x"09",x"71",x"d4",x"d8",x"d8",x"d8",x"b4",x"6c",x"b0",x"d8",x"d8",x"d8",x"f8",x"b5",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"b5",x"8d",x"91",x"99",x"78",x"55",x"75",x"b8",x"75",x"0e",x"11",x"51",x"50",x"51",x"55",x"0d",x"0d",x"0d",x"0d",x"55",x"b9",x"99",x"75",x"70",x"99",x"75",x"78",x"75",x"31",x"12",x"15",x"16",x"16",x"16",x"11",x"0d",x"16",x"12",x"12",x"2d",x"2c",x"2c",x"2c",x"0d",x"12",x"11",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"0d",x"11",x"11",x"11",x"15",x"11",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"11"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"0d",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"32",x"2e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2e",x"2d",x"2d",x"4d",x"4d",x"2d",x"49",x"49",x"4d",x"49",x"49",x"2d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"0e",x"75",x"98",x"55",x"12",x"16",x"16",x"99",x"98",x"98",x"79",x"75",x"55",x"55",x"55",x"55",x"15",x"16",x"16",x"16",x"16",x"55",x"79",x"98",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"71",x"90",x"90",x"90",x"d8",x"fc",x"d8",x"94",x"90",x"71",x"70",x"6c",x"70",x"94",x"b4",x"b4",x"b8",x"d4",x"d8",x"b4",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"8d",x"d5",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"49",x"b1",x"b5",x"d1",x"92",x"13",x"12",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"b4",x"b4",x"b4",x"b4",x"90",x"6c",x"90",x"d4",x"d8",x"d8",x"f8",x"b5",x"2e",x"0d",x"0e",x"0d",x"0d",x"0d",x"0e",x"0d",x"0e",x"0e",x"0d",x"0e",x"0d",x"0d",x"0e",x"12",x"b1",x"6d",x"91",x"98",x"98",x"55",x"55",x"b8",x"95",x"12",x"11",x"55",x"54",x"55",x"55",x"0d",x"11",x"0d",x"11",x"75",x"b9",x"99",x"75",x"71",x"99",x"75",x"75",x"75",x"55",x"12",x"11",x"12",x"11",x"16",x"11",x"0d",x"16",x"15",x"12",x"0d",x"28",x"28",x"0d",x"0d",x"11",x"11",x"11",x"12",x"16",x"11",x"0d",x"0d",x"11",x"0d",x"12",x"11",x"15",x"15",x"15",x"16",x"16",x"16",x"12",x"11",x"0d",x"0d",x"09",x"05"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"0d",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"0d",x"11",x"12",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2d",x"2d",x"29",x"29",x"29",x"2d",x"49",x"49",x"2d",x"29",x"29",x"2d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0e",x"55",x"98",x"75",x"12",x"16",x"16",x"99",x"98",x"98",x"99",x"75",x"55",x"55",x"75",x"55",x"15",x"16",x"16",x"12",x"0d",x"75",x"75",x"99",x"2d",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0e",x"0a",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"4d",x"90",x"90",x"90",x"94",x"d8",x"fd",x"d8",x"b4",x"70",x"70",x"70",x"70",x"70",x"90",x"90",x"94",x"b4",x"b4",x"95",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"91",x"b1",x"d1",x"b1",x"b1",x"b1",x"b1",x"71",x"b1",x"b5",x"d1",x"72",x"12",x"12",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0e",x"12",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"4d",x"90",x"b4",x"90",x"90",x"6c",x"90",x"b4",x"b4",x"d4",x"f8",x"b5",x"0e",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"12",x"11",x"12",x"11",x"11",x"12",x"12",x"91",x"6d",x"91",x"99",x"98",x"55",x"51",x"b8",x"99",x"12",x"31",x"55",x"50",x"50",x"55",x"0d",x"0d",x"0d",x"31",x"75",x"b9",x"99",x"75",x"71",x"99",x"75",x"75",x"75",x"55",x"12",x"12",x"12",x"15",x"16",x"11",x"0d",x"16",x"12",x"12",x"09",x"08",x"08",x"0d",x"11",x"11",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"16",x"16",x"16",x"16",x"11",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"05",x"05"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"0d",x"0d",x"12",x"32",x"52",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"2d",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"31",x"75",x"99",x"35",x"16",x"16",x"75",x"98",x"98",x"98",x"75",x"55",x"55",x"54",x"55",x"15",x"12",x"11",x"09",x"09",x"75",x"79",x"79",x"2d",x"09",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"2e",x"4d",x"4e",x"2e",x"2e",x"0e",x"2d",x"71",x"90",x"90",x"70",x"b4",x"d8",x"d8",x"d9",x"b5",x"70",x"70",x"70",x"70",x"70",x"70",x"70",x"91",x"90",x"91",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4e",x"91",x"b1",x"b1",x"b5",x"b5",x"b5",x"91",x"b1",x"b5",x"b1",x"72",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"0e",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"91",x"90",x"90",x"70",x"6c",x"90",x"90",x"94",x"b4",x"d4",x"95",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"12",x"11",x"12",x"12",x"12",x"12",x"12",x"91",x"6d",x"91",x"95",x"99",x"55",x"51",x"b9",x"98",x"12",x"31",x"55",x"54",x"51",x"55",x"0d",x"11",x"11",x"31",x"95",x"b9",x"99",x"75",x"70",x"99",x"75",x"75",x"74",x"55",x"12",x"12",x"12",x"16",x"16",x"11",x"0d",x"11",x"12",x"11",x"08",x"04",x"08",x"0d",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"11",x"12",x"12",x"16",x"11",x"12",x"12",x"11",x"0d",x"0d",x"09",x"05",x"05",x"05",x"05",x"05",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"11",x"11",x"11",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"12",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"32",x"2e",x"2e",x"2e",x"4e",x"4e",x"2d",x"4d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"49",x"2d",x"49",x"45",x"29",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"55",x"98",x"75",x"16",x"16",x"75",x"98",x"98",x"99",x"74",x"55",x"55",x"55",x"55",x"0d",x"09",x"09",x"09",x"09",x"78",x"78",x"75",x"2d",x"09",x"09",x"09",x"09",x"0d",x"0a",x"0e",x"71",x"d4",x"d8",x"d8",x"b5",x"91",x"70",x"70",x"90",x"90",x"91",x"70",x"b5",x"d4",x"d8",x"d8",x"b4",x"90",x"70",x"70",x"70",x"70",x"70",x"70",x"90",x"95",x"2d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"8d",x"b1",x"b1",x"b1",x"6d",x"b1",x"b1",x"8d",x"4e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"1a",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0e",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"6d",x"90",x"70",x"70",x"6c",x"70",x"90",x"90",x"b4",x"b4",x"71",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"12",x"12",x"12",x"12",x"71",x"6d",x"91",x"95",x"99",x"75",x"31",x"99",x"b8",x"36",x"35",x"55",x"55",x"55",x"55",x"12",x"16",x"12",x"35",x"99",x"b9",x"99",x"51",x"50",x"99",x"75",x"75",x"74",x"55",x"11",x"12",x"16",x"16",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"08",x"04",x"0d",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"0d",x"09",x"09",x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"11",x"11",x"0d",x"0d",x"11",x"11",x"11",x"11",x"0e",x"32",x"32",x"2e",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"49",x"29",x"29",x"29",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"55",x"98",x"79",x"16",x"16",x"55",x"98",x"98",x"98",x"98",x"75",x"55",x"55",x"55",x"0d",x"09",x"09",x"09",x"2d",x"78",x"78",x"55",x"0d",x"09",x"09",x"09",x"09",x"0e",x"0a",x"71",x"d8",x"d8",x"d8",x"d8",x"d4",x"b0",x"90",x"90",x"90",x"70",x"70",x"70",x"90",x"b4",x"d8",x"d8",x"b4",x"90",x"90",x"70",x"70",x"70",x"70",x"70",x"90",x"91",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"8d",x"8d",x"6d",x"49",x"8d",x"8d",x"6d",x"2e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"17",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"12",x"0e",x"12",x"13",x"13",x"13",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"4d",x"70",x"70",x"6c",x"6c",x"70",x"90",x"b0",x"90",x"4d",x"2d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"12",x"71",x"6d",x"91",x"95",x"99",x"75",x"31",x"79",x"98",x"56",x"55",x"55",x"55",x"55",x"55",x"16",x"16",x"16",x"55",x"95",x"99",x"99",x"51",x"71",x"99",x"75",x"75",x"74",x"75",x"35",x"12",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"11",x"08",x"08",x"08",x"11",x"16",x"16",x"16",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"0d",x"12",x"32",x"32",x"32",x"2e",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2d",x"2d",x"2d",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"16",x"16",x"35",x"75",x"75",x"35",x"16",x"35",x"75",x"75",x"95",x"95",x"75",x"55",x"74",x"55",x"09",x"09",x"09",x"09",x"2d",x"79",x"78",x"51",x"09",x"09",x"09",x"09",x"09",x"0e",x"2e",x"b4",x"f8",x"d8",x"b4",x"d4",x"d4",x"b4",x"b4",x"90",x"90",x"70",x"70",x"90",x"90",x"90",x"b4",x"b4",x"b4",x"94",x"90",x"70",x"70",x"70",x"90",x"90",x"94",x"95",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4d",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"2e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"12",x"12",x"0e",x"12",x"13",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"11",x"11",x"12",x"11",x"31",x"31",x"31",x"31",x"11",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"4d",x"70",x"70",x"6c",x"70",x"70",x"90",x"90",x"4d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"12",x"12",x"12",x"12",x"71",x"6d",x"91",x"95",x"99",x"75",x"31",x"75",x"98",x"55",x"55",x"54",x"55",x"55",x"55",x"16",x"16",x"16",x"55",x"95",x"99",x"99",x"51",x"71",x"99",x"75",x"75",x"75",x"75",x"35",x"12",x"11",x"0d",x"11",x"0d",x"0d",x"11",x"11",x"08",x"08",x"0d",x"11",x"16",x"11",x"11",x"0d",x"0d",x"0d",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"0e",x"2e",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"2d",x"2d",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"0d",x"11",x"11",x"11",x"11",x"0d",x"11",x"16",x"16",x"16",x"16",x"11",x"12",x"11",x"11",x"11",x"16",x"15",x"32",x"32",x"4e",x"4d",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"4e",x"51",x"51",x"55",x"54",x"74",x"09",x"09",x"09",x"09",x"51",x"79",x"78",x"51",x"09",x"09",x"09",x"09",x"0e",x"0a",x"51",x"b4",x"d8",x"d8",x"d4",x"d4",x"d8",x"b4",x"94",x"90",x"70",x"70",x"90",x"90",x"90",x"71",x"91",x"b4",x"b4",x"94",x"91",x"70",x"70",x"90",x"94",x"94",x"b4",x"b4",x"4e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4d",x"6d",x"6d",x"49",x"4d",x"6d",x"6d",x"2e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"13",x"17",x"17",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"13",x"13",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"1a",x"1a",x"1a",x"1a",x"1a",x"1a",x"1a",x"1a",x"1a",x"1a",x"16",x"1a",x"16",x"16",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"32",x"51",x"55",x"75",x"75",x"74",x"74",x"70",x"70",x"70",x"70",x"70",x"51",x"31",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"09",x"09",x"0d",x"09",x"09",x"4d",x"70",x"70",x"6c",x"70",x"70",x"90",x"2d",x"09",x"09",x"09",x"0d",x"0d",x"12",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"71",x"6d",x"8d",x"95",x"99",x"74",x"51",x"75",x"98",x"75",x"55",x"55",x"54",x"55",x"55",x"16",x"16",x"12",x"55",x"75",x"99",x"99",x"51",x"50",x"99",x"75",x"55",x"75",x"75",x"55",x"12",x"16",x"16",x"16",x"11",x"11",x"11",x"09",x"08",x"08",x"0d",x"0d",x"09",x"09",x"05",x"05",x"09",x"09",x"09",x"05",x"05",x"09",x"09",x"05",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"09",x"0d",x"11",x"11",x"11",x"11",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"31",x"2d",x"4d",x"4d",x"4e",x"2d",x"2a",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"51",x"51",x"51",x"2d",x"09",x"09",x"09",x"55",x"75",x"78",x"2d",x"09",x"09",x"09",x"09",x"0a",x"0a",x"71",x"d8",x"d8",x"d8",x"d8",x"d4",x"d8",x"94",x"70",x"70",x"90",x"90",x"70",x"90",x"51",x"2e",x"71",x"b4",x"d8",x"b4",x"94",x"6c",x"70",x"90",x"94",x"b4",x"b8",x"d8",x"95",x"52",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"4d",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"55",x"75",x"75",x"75",x"95",x"95",x"94",x"94",x"94",x"94",x"70",x"70",x"70",x"70",x"70",x"51",x"31",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"4d",x"90",x"90",x"70",x"6c",x"70",x"90",x"90",x"2d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"71",x"6d",x"8d",x"91",x"99",x"78",x"55",x"51",x"99",x"75",x"75",x"55",x"55",x"75",x"55",x"16",x"16",x"12",x"55",x"75",x"95",x"99",x"50",x"50",x"95",x"75",x"55",x"55",x"75",x"55",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"08",x"08",x"08",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"11",x"0d",x"11",x"11",x"0d",x"0d",x"11",x"11",x"2e",x"32",x"32",x"32",x"2e",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"49",x"49",x"25",x"25",x"29",x"0d",x"11",x"11",x"11",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"4d",x"49",x"4d",x"4d",x"4e",x"4d",x"4d",x"4e",x"4e",x"4d",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"0d",x"09",x"09",x"75",x"74",x"79",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"71",x"b4",x"d8",x"d8",x"d8",x"d4",x"b4",x"90",x"6c",x"70",x"94",x"b4",x"90",x"71",x"0e",x"0e",x"95",x"d8",x"d8",x"d4",x"94",x"6c",x"70",x"94",x"b4",x"b8",x"b8",x"d8",x"d8",x"95",x"4e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"4e",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"17",x"13",x"13",x"13",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0e",x"0d",x"0e",x"0d",x"0d",x"0e",x"0d",x"11",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"36",x"55",x"95",x"95",x"b4",x"94",x"94",x"94",x"95",x"75",x"70",x"71",x"75",x"71",x"70",x"70",x"71",x"71",x"70",x"50",x"2d",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"2d",x"4d",x"94",x"b4",x"94",x"90",x"70",x"70",x"74",x"71",x"51",x"31",x"31",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"71",x"91",x"6d",x"91",x"95",x"78",x"55",x"51",x"99",x"75",x"75",x"55",x"55",x"75",x"59",x"16",x"16",x"12",x"51",x"74",x"75",x"99",x"70",x"50",x"75",x"75",x"54",x"55",x"75",x"75",x"0d",x"0d",x"09",x"09",x"09",x"08",x"09",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"2d",x"2d",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"11",x"0d",x"0d",x"11",x"0d",x"0d",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"2d",x"2d",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"49",x"29",x"29",x"29",x"29",x"25",x"29",x"11",x"11",x"11",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"49",x"49",x"4e",x"4d",x"4e",x"4e",x"4e",x"4e",x"2e",x"29",x"4d",x"4e",x"4e",x"2e",x"2e",x"4e",x"2e",x"2e",x"2e",x"2e",x"32",x"2e",x"2e",x"55",x"74",x"78",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"4d",x"b4",x"d8",x"d8",x"d9",x"b4",x"70",x"94",x"b4",x"b4",x"94",x"b4",x"91",x"2e",x"0e",x"95",x"d4",x"b4",x"d4",x"d8",x"b4",x"6c",x"70",x"94",x"b4",x"d4",x"b4",x"b8",x"b4",x"b8",x"b4",x"52",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"4d",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"09",x"09",x"0a",x"0a",x"0a",x"0a",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"12",x"16",x"16",x"16",x"36",x"75",x"95",x"98",x"94",x"94",x"94",x"95",x"94",x"94",x"95",x"70",x"70",x"71",x"75",x"74",x"71",x"70",x"71",x"71",x"70",x"70",x"2c",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"51",x"b5",x"d4",x"b8",x"b8",x"95",x"95",x"75",x"75",x"55",x"51",x"51",x"51",x"74",x"74",x"75",x"75",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"51",x"91",x"6d",x"8d",x"95",x"99",x"55",x"31",x"99",x"75",x"75",x"55",x"55",x"75",x"59",x"16",x"16",x"12",x"31",x"70",x"75",x"75",x"75",x"51",x"75",x"55",x"54",x"55",x"55",x"51",x"09",x"05",x"09",x"09",x"09",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"05",x"2d",x"50",x"2d",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"0d",x"2d",x"2e",x"32",x"32",x"2e",x"32",x"32",x"2e",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"2d",x"2d",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"49",x"49",x"29",x"24",x"0d",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"11",x"2d",x"49",x"49",x"2d",x"4d",x"4d",x"2d",x"2d",x"4d",x"29",x"2d",x"4e",x"2e",x"2e",x"4e",x"4e",x"4e",x"2e",x"2e",x"2e",x"4e",x"52",x"32",x"52",x"52",x"51",x"75",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"90",x"d8",x"d8",x"d9",x"94",x"90",x"b4",x"d8",x"b4",x"b4",x"b4",x"91",x"0e",x"71",x"d4",x"d8",x"b8",x"b8",x"b8",x"b4",x"70",x"70",x"94",x"b4",x"b8",x"b4",x"b4",x"b4",x"b8",x"d8",x"71",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"09",x"09",x"0a",x"09",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"16",x"1a",x"36",x"55",x"75",x"95",x"b8",x"b8",x"94",x"95",x"95",x"94",x"95",x"95",x"95",x"74",x"71",x"71",x"50",x"50",x"71",x"70",x"50",x"50",x"50",x"4c",x"2c",x"0d",x"12",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"0d",x"11",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"51",x"b5",x"d8",x"b8",x"94",x"75",x"75",x"55",x"75",x"55",x"75",x"75",x"94",x"94",x"94",x"98",x"95",x"95",x"55",x"31",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"51",x"91",x"6d",x"8d",x"95",x"99",x"75",x"31",x"99",x"75",x"55",x"55",x"55",x"75",x"55",x"12",x"12",x"0e",x"31",x"50",x"75",x"75",x"75",x"4d",x"75",x"55",x"55",x"51",x"75",x"51",x"29",x"05",x"09",x"09",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"2c",x"50",x"2d",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"11",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"2d",x"2e",x"32",x"32",x"2e",x"32",x"32",x"2e",x"32",x"32",x"2e",x"2e",x"2e",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"2d",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"49",x"4d",x"4d",x"4d",x"24",x"29",x"11",x"16",x"16",x"16",x"16",x"16",x"11",x"0d",x"09",x"29",x"29",x"4d",x"29",x"29",x"49",x"29",x"29",x"29",x"29",x"4e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2e",x"2d",x"2d",x"2d",x"2e",x"32",x"32",x"2e",x"2e",x"32",x"52",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"71",x"b4",x"b8",x"b4",x"94",x"d4",x"d8",x"d8",x"d8",x"b4",x"b4",x"71",x"0e",x"b4",x"d8",x"b8",x"b8",x"b8",x"b8",x"b4",x"70",x"6c",x"94",x"b4",x"b8",x"b8",x"b4",x"b8",x"b4",x"d8",x"b5",x"4d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"6d",x"8d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"8d",x"6d",x"2e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"16",x"3a",x"79",x"b8",x"b8",x"b8",x"98",x"94",x"94",x"95",x"95",x"94",x"95",x"95",x"75",x"75",x"75",x"70",x"4c",x"4c",x"50",x"51",x"50",x"50",x"50",x"4c",x"2c",x"2d",x"12",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"2d",x"95",x"f8",x"94",x"75",x"75",x"51",x"50",x"50",x"50",x"75",x"94",x"98",x"b8",x"b8",x"b8",x"b8",x"98",x"95",x"94",x"75",x"51",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"52",x"91",x"6d",x"8d",x"91",x"99",x"75",x"31",x"99",x"55",x"55",x"55",x"55",x"74",x"71",x"09",x"09",x"09",x"2d",x"50",x"75",x"55",x"50",x"2c",x"51",x"55",x"55",x"51",x"54",x"54",x"2d",x"09",x"09",x"09",x"08",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"31",x"51",x"50",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"2d",x"2e",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2d",x"29",x"29",x"29",x"49",x"29",x"29",x"49",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"29",x"24",x"2d",x"16",x"16",x"11",x"0d",x"0d",x"09",x"09",x"09",x"29",x"49",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"49",x"29",x"29",x"29",x"2d",x"2d",x"2d",x"2d",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"2e",x"09",x"09",x"09",x"0d",x"09",x"09",x"71",x"b4",x"94",x"90",x"b8",x"d8",x"d8",x"b4",x"b4",x"d8",x"b4",x"94",x"2e",x"d4",x"d4",x"b4",x"b4",x"b4",x"b8",x"b4",x"70",x"6c",x"90",x"b4",x"b8",x"b4",x"b4",x"b4",x"b8",x"d8",x"b5",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"b1",x"8d",x"8d",x"6d",x"6d",x"6d",x"6d",x"29",x"6d",x"8d",x"4d",x"2e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"55",x"99",x"b8",x"b8",x"b8",x"b8",x"98",x"94",x"94",x"75",x"70",x"70",x"70",x"70",x"70",x"71",x"71",x"71",x"70",x"50",x"2c",x"51",x"51",x"50",x"50",x"2c",x"2c",x"0d",x"12",x"12",x"11",x"12",x"12",x"11",x"11",x"11",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0e",x"51",x"95",x"94",x"75",x"50",x"51",x"75",x"99",x"98",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"d8",x"dd",x"b9",x"b9",x"95",x"55",x"11",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"56",x"91",x"6d",x"6d",x"91",x"b9",x"75",x"30",x"75",x"75",x"75",x"55",x"54",x"75",x"55",x"09",x"09",x"09",x"2d",x"51",x"51",x"51",x"50",x"2c",x"50",x"55",x"51",x"51",x"51",x"51",x"2d",x"09",x"09",x"09",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"2d",x"31",x"30",x"51",x"50",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"2d",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2d",x"2d",x"2d",x"4d",x"4d",x"4d",x"29",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"24",x"29",x"11",x"11",x"0d",x"09",x"09",x"09",x"09",x"09",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2d",x"2d",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"0d",x"09",x"0d",x"0d",x"09",x"71",x"94",x"90",x"70",x"d8",x"d9",x"d8",x"d8",x"d8",x"d8",x"d8",x"b4",x"71",x"d8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b4",x"70",x"6c",x"90",x"b4",x"b8",x"b8",x"b8",x"b8",x"b8",x"d8",x"b5",x"51",x"0a",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"b1",x"8d",x"8d",x"8d",x"8d",x"8d",x"6d",x"49",x"49",x"8d",x"8d",x"4e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0d",x"0d",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"51",x"95",x"b8",x"b8",x"b8",x"b8",x"98",x"98",x"94",x"94",x"94",x"74",x"71",x"71",x"70",x"70",x"50",x"4c",x"51",x"50",x"50",x"4c",x"4c",x"50",x"50",x"4c",x"2c",x"2c",x"0d",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"51",x"74",x"75",x"74",x"74",x"74",x"99",x"b8",x"b8",x"b8",x"d8",x"b8",x"b8",x"b8",x"b4",x"95",x"75",x"75",x"95",x"b9",x"b9",x"b9",x"99",x"75",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"32",x"91",x"91",x"6d",x"91",x"b5",x"75",x"30",x"75",x"75",x"75",x"55",x"55",x"75",x"55",x"09",x"09",x"09",x"2d",x"51",x"51",x"55",x"51",x"2c",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"05",x"05",x"05",x"08",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"0d",x"2d",x"2d",x"30",x"50",x"2c",x"51",x"51",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"12",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"0d",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"29",x"2e",x"32",x"32",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2d",x"2d",x"4e",x"4e",x"4e",x"4d",x"2d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"52",x"29",x"25",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"25",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2d",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"52",x"32",x"32",x"32",x"2e",x"09",x"0d",x"0d",x"0a",x"4d",x"90",x"70",x"70",x"d8",x"d9",x"d8",x"d9",x"d8",x"d8",x"d8",x"d4",x"95",x"b8",x"b8",x"b8",x"b8",x"b8",x"d8",x"b4",x"70",x"4c",x"90",x"b4",x"b8",x"d8",x"d8",x"b9",x"d8",x"d8",x"91",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"b1",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"29",x"6d",x"ad",x"6d",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"51",x"b9",x"b8",x"b8",x"b8",x"98",x"98",x"98",x"98",x"94",x"94",x"94",x"95",x"95",x"95",x"71",x"70",x"50",x"4c",x"4c",x"2c",x"4c",x"50",x"2c",x"4c",x"50",x"4c",x"2c",x"2d",x"11",x"12",x"11",x"12",x"11",x"11",x"11",x"12",x"0e",x"11",x"11",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"51",x"75",x"54",x"75",x"98",x"b8",x"b8",x"b8",x"94",x"90",x"b4",x"d8",x"d4",x"b4",x"b4",x"d4",x"51",x"0e",x"0e",x"32",x"76",x"99",x"b9",x"b9",x"b9",x"75",x"11",x"16",x"16",x"12",x"12",x"12",x"11",x"0e",x"0e",x"91",x"91",x"6d",x"91",x"b5",x"79",x"31",x"55",x"75",x"75",x"55",x"55",x"75",x"75",x"09",x"0d",x"09",x"2d",x"51",x"51",x"55",x"51",x"2c",x"51",x"50",x"50",x"71",x"71",x"71",x"71",x"09",x"05",x"05",x"08",x"08",x"09",x"09",x"09",x"09",x"08",x"09",x"09",x"09",x"0d",x"2d",x"2d",x"2d",x"31",x"50",x"50",x"30",x"2c",x"2c",x"75",x"51",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"12",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"29",x"2d",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"2d",x"4e",x"2e",x"2e",x"4e",x"4e",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"09",x"24",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"45",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2d",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"09",x"0d",x"09",x"4d",x"90",x"90",x"70",x"b4",x"b8",x"d8",x"d9",x"d9",x"d8",x"d8",x"d8",x"95",x"d8",x"d9",x"d9",x"d9",x"d9",x"d9",x"b8",x"90",x"4c",x"70",x"b4",x"b8",x"b8",x"b8",x"b4",x"94",x"94",x"4d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"b1",x"91",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"49",x"69",x"8d",x"8d",x"4e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"51",x"99",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"99",x"95",x"95",x"94",x"94",x"94",x"75",x"71",x"71",x"70",x"70",x"70",x"50",x"50",x"4c",x"2c",x"2c",x"2c",x"2c",x"29",x"11",x"12",x"12",x"12",x"16",x"12",x"12",x"0d",x"0d",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"36",x"36",x"36",x"75",x"75",x"94",x"98",x"b8",x"b8",x"d8",x"d8",x"b4",x"70",x"70",x"b4",x"d8",x"d8",x"d8",x"d8",x"d8",x"75",x"12",x"12",x"16",x"16",x"36",x"55",x"75",x"94",x"99",x"75",x"32",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"8d",x"91",x"6d",x"91",x"b5",x"75",x"51",x"51",x"75",x"75",x"75",x"55",x"74",x"75",x"09",x"0e",x"0e",x"0d",x"31",x"51",x"51",x"70",x"70",x"94",x"94",x"b4",x"b8",x"b8",x"b8",x"b4",x"71",x"4d",x"50",x"28",x"04",x"05",x"09",x"08",x"2c",x"2c",x"2c",x"2c",x"2d",x"2c",x"2d",x"2c",x"2c",x"30",x"30",x"50",x"30",x"08",x"50",x"74",x"2d",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"2d",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"2e",x"2e",x"4e",x"2e",x"2e",x"2e",x"4e",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"09",x"04",x"24",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2d",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"52",x"32",x"0d",x"0d",x"09",x"4d",x"90",x"70",x"70",x"94",x"b4",x"d8",x"d9",x"d9",x"d8",x"d8",x"d9",x"95",x"b5",x"d8",x"d9",x"d9",x"d9",x"d9",x"b8",x"94",x"4c",x"70",x"94",x"b4",x"b4",x"94",x"94",x"94",x"71",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"91",x"b1",x"91",x"8d",x"8d",x"8d",x"8d",x"8d",x"69",x"49",x"6d",x"ad",x"6d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0a",x"0a",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"31",x"99",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"99",x"99",x"94",x"94",x"94",x"94",x"75",x"70",x"71",x"70",x"70",x"50",x"50",x"4d",x"4c",x"2c",x"2c",x"2c",x"2c",x"2d",x"0d",x"0d",x"12",x"16",x"16",x"12",x"12",x"11",x"11",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"32",x"35",x"55",x"55",x"75",x"99",x"94",x"94",x"b8",x"b8",x"b8",x"b4",x"d4",x"90",x"6c",x"70",x"b4",x"d8",x"d8",x"d8",x"d8",x"d8",x"75",x"12",x"11",x"11",x"16",x"12",x"11",x"31",x"54",x"74",x"94",x"75",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"6d",x"91",x"6d",x"8d",x"b5",x"95",x"55",x"31",x"55",x"75",x"75",x"55",x"74",x"75",x"0a",x"0e",x"0e",x"0e",x"2d",x"51",x"71",x"94",x"94",x"94",x"94",x"94",x"b4",x"d8",x"d8",x"d8",x"d8",x"b4",x"94",x"50",x"2c",x"29",x"08",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"08",x"75",x"50",x"2d",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"09",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"2d",x"32",x"2e",x"2e",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2d",x"29",x"4d",x"2d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"09",x"05",x"24",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"4e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"09",x"29",x"6d",x"70",x"70",x"90",x"94",x"94",x"b4",x"b8",x"d8",x"d8",x"d8",x"d9",x"95",x"75",x"b8",x"d8",x"d8",x"d9",x"b8",x"b4",x"90",x"4c",x"70",x"90",x"91",x"90",x"90",x"90",x"90",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"52",x"b1",x"b5",x"b1",x"91",x"91",x"91",x"91",x"8d",x"49",x"6d",x"ad",x"6d",x"2e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"95",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"98",x"98",x"98",x"98",x"94",x"95",x"95",x"70",x"70",x"70",x"50",x"4c",x"4c",x"4c",x"4c",x"4c",x"2c",x"2c",x"2c",x"2c",x"2c",x"28",x"28",x"31",x"12",x"16",x"16",x"16",x"11",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"55",x"75",x"75",x"75",x"95",x"95",x"95",x"b8",x"98",x"94",x"91",x"b0",x"b4",x"90",x"70",x"6c",x"90",x"b4",x"d4",x"d8",x"d8",x"b4",x"d8",x"71",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"2d",x"51",x"55",x"75",x"99",x"51",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"6d",x"91",x"8d",x"8d",x"b1",x"95",x"55",x"31",x"55",x"79",x"75",x"55",x"75",x"79",x"0e",x"0e",x"0e",x"0e",x"2d",x"75",x"b4",x"b8",x"94",x"70",x"70",x"4c",x"6c",x"90",x"b4",x"fc",x"fc",x"d8",x"b4",x"94",x"b8",x"70",x"08",x"08",x"08",x"28",x"28",x"2c",x"2c",x"28",x"2c",x"2c",x"2c",x"2c",x"2c",x"08",x"08",x"2c",x"75",x"51",x"0d",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05"),
(x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"2d",x"4d",x"6d",x"8d",x"8d",x"8d",x"6d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0e",x"0d",x"0d",x"0e",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"2d",x"2d",x"32",x"32",x"2e",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"2d",x"4e",x"2d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"2d",x"09",x"05",x"24",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2d",x"2d",x"2d",x"2d",x"2d",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"29",x"4d",x"70",x"70",x"6c",x"70",x"91",x"94",x"94",x"b4",x"b4",x"d8",x"d8",x"d8",x"95",x"2e",x"75",x"b4",x"b4",x"b4",x"94",x"94",x"90",x"6c",x"6c",x"70",x"70",x"70",x"94",x"90",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"91",x"b1",x"b1",x"b5",x"b5",x"b5",x"91",x"71",x"91",x"8d",x"6d",x"2e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"b8",x"b8",x"b8",x"b8",x"b9",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"94",x"94",x"74",x"75",x"75",x"71",x"50",x"50",x"51",x"51",x"50",x"50",x"51",x"4c",x"2c",x"2c",x"2c",x"50",x"4c",x"4c",x"2c",x"2c",x"2d",x"11",x"16",x"16",x"15",x"16",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"51",x"75",x"71",x"75",x"75",x"95",x"b9",x"98",x"74",x"70",x"71",x"75",x"90",x"90",x"90",x"6c",x"6c",x"70",x"94",x"b4",x"b4",x"d8",x"d8",x"d8",x"6d",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"2d",x"55",x"55",x"75",x"99",x"4d",x"0a",x"09",x"0d",x"0d",x"09",x"4d",x"91",x"91",x"8d",x"91",x"b5",x"54",x"30",x"55",x"75",x"74",x"55",x"75",x"75",x"0e",x"0e",x"0d",x"0e",x"51",x"95",x"94",x"70",x"71",x"4c",x"4c",x"4c",x"4c",x"4c",x"50",x"70",x"94",x"dc",x"dc",x"b8",x"b4",x"94",x"70",x"28",x"08",x"28",x"2c",x"2c",x"28",x"2c",x"2c",x"2c",x"2c",x"28",x"08",x"08",x"28",x"75",x"75",x"31",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"05",x"05",x"05"),
(x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"4d",x"8d",x"ad",x"cc",x"cc",x"cc",x"cc",x"cc",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"6d",x"6d",x"6d",x"4d",x"4d",x"2d",x"2d",x"0d",x"0d",x"2d",x"4d",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"2d",x"2e",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4e",x"09",x"09",x"09",x"24",x"25",x"09",x"09",x"09",x"09",x"0d",x"09",x"29",x"29",x"49",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2d",x"2d",x"2d",x"2e",x"2d",x"2d",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"29",x"70",x"70",x"70",x"6c",x"70",x"91",x"90",x"90",x"94",x"b4",x"b4",x"d8",x"b4",x"51",x"0a",x"2e",x"71",x"94",x"94",x"94",x"90",x"70",x"6c",x"4c",x"6c",x"70",x"70",x"90",x"94",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4d",x"6d",x"8d",x"91",x"91",x"91",x"b1",x"91",x"71",x"91",x"8d",x"6d",x"2e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"32",x"95",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"94",x"94",x"94",x"94",x"94",x"74",x"74",x"74",x"74",x"70",x"50",x"51",x"71",x"50",x"51",x"50",x"4c",x"4c",x"4c",x"4c",x"50",x"50",x"50",x"2c",x"2c",x"28",x"2d",x"11",x"12",x"11",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"31",x"71",x"75",x"51",x"75",x"75",x"95",x"99",x"94",x"50",x"50",x"51",x"75",x"90",x"70",x"70",x"6c",x"6c",x"6c",x"90",x"94",x"b4",x"b4",x"b4",x"b4",x"4d",x"05",x"09",x"05",x"09",x"0e",x"0d",x"0a",x"0d",x"31",x"55",x"55",x"78",x"75",x"2d",x"09",x"09",x"0d",x"09",x"4d",x"91",x"b1",x"8d",x"8d",x"b5",x"74",x"2c",x"55",x"75",x"74",x"55",x"75",x"75",x"0e",x"0e",x"0d",x"0e",x"71",x"94",x"70",x"4c",x"51",x"4c",x"4c",x"4c",x"4c",x"2c",x"2c",x"2d",x"4c",x"94",x"dc",x"d8",x"b4",x"b4",x"94",x"6c",x"28",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"28",x"08",x"08",x"28",x"51",x"75",x"50",x"2d",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"05",x"05",x"05",x"05"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"4d",x"ac",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"6d",x"11",x"0d",x"0d",x"0d",x"0d",x"89",x"e8",x"e8",x"e8",x"e8",x"ec",x"cc",x"ad",x"11",x"6d",x"cc",x"cc",x"8d",x"4d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"29",x"2d",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"2e",x"2e",x"4e",x"4e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4e",x"2e",x"09",x"09",x"09",x"24",x"25",x"09",x"09",x"09",x"09",x"0d",x"29",x"49",x"29",x"29",x"49",x"29",x"29",x"29",x"29",x"29",x"49",x"29",x"29",x"29",x"29",x"4e",x"2e",x"2e",x"2e",x"2e",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"29",x"4d",x"70",x"6c",x"6c",x"70",x"70",x"70",x"70",x"90",x"90",x"94",x"94",x"71",x"09",x"09",x"09",x"0d",x"71",x"94",x"90",x"90",x"70",x"6c",x"4c",x"6c",x"70",x"70",x"70",x"94",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"29",x"69",x"8d",x"8d",x"6d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"11",x"11",x"11",x"12",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"99",x"94",x"94",x"74",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"71",x"71",x"70",x"50",x"71",x"2c",x"2c",x"51",x"4c",x"4c",x"50",x"51",x"4c",x"50",x"50",x"4c",x"28",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"2d",x"31",x"51",x"55",x"51",x"75",x"95",x"95",x"75",x"50",x"50",x"70",x"74",x"74",x"91",x"70",x"70",x"6c",x"6c",x"70",x"70",x"70",x"90",x"90",x"94",x"91",x"29",x"05",x"09",x"09",x"09",x"0e",x"0e",x"0e",x"0e",x"11",x"74",x"50",x"51",x"74",x"51",x"0d",x"09",x"0d",x"09",x"2d",x"91",x"b5",x"8d",x"8d",x"b5",x"75",x"2c",x"55",x"75",x"74",x"50",x"75",x"79",x"2e",x"0e",x"0e",x"71",x"70",x"70",x"50",x"71",x"71",x"70",x"4c",x"2d",x"30",x"2d",x"2d",x"2d",x"08",x"04",x"94",x"fc",x"dc",x"b4",x"71",x"b4",x"50",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"0c",x"2c",x"71",x"75",x"75",x"50",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"09"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"12",x"12",x"11",x"11",x"11",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"cc",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"4d",x"0e",x"0e",x"0d",x"0d",x"0e",x"89",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"6d",x"89",x"c8",x"e8",x"cc",x"cc",x"8c",x"6d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"29",x"2e",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"2e",x"2e",x"4e",x"4e",x"4e",x"4d",x"4d",x"4d",x"4d",x"4e",x"52",x"2d",x"09",x"09",x"09",x"09",x"24",x"24",x"09",x"09",x"09",x"09",x"2d",x"49",x"49",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2d",x"2d",x"2e",x"2e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"29",x"71",x"70",x"6c",x"6c",x"70",x"70",x"70",x"70",x"71",x"4d",x"2d",x"2d",x"29",x"0d",x"0d",x"12",x"16",x"16",x"55",x"94",x"70",x"70",x"6c",x"4c",x"4c",x"70",x"70",x"70",x"90",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"29",x"6d",x"6d",x"6d",x"4e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2d",x"75",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"98",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"95",x"75",x"70",x"70",x"50",x"4c",x"4c",x"50",x"50",x"4c",x"2c",x"50",x"4d",x"51",x"50",x"50",x"50",x"2c",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0e",x"2d",x"31",x"51",x"51",x"75",x"75",x"75",x"51",x"51",x"51",x"51",x"71",x"75",x"74",x"70",x"90",x"70",x"6c",x"6c",x"70",x"70",x"6c",x"90",x"90",x"94",x"95",x"75",x"51",x"09",x"05",x"09",x"0e",x"0e",x"0e",x"0e",x"0d",x"51",x"74",x"55",x"50",x"75",x"2d",x"0a",x"0d",x"09",x"09",x"91",x"b5",x"91",x"6d",x"b5",x"95",x"30",x"55",x"75",x"75",x"51",x"54",x"75",x"31",x"0e",x"51",x"71",x"70",x"70",x"70",x"70",x"71",x"50",x"2d",x"2d",x"2c",x"2c",x"2c",x"2c",x"08",x"04",x"28",x"94",x"dc",x"d8",x"94",x"70",x"94",x"70",x"28",x"08",x"28",x"2c",x"2c",x"2c",x"50",x"51",x"75",x"75",x"75",x"50",x"2d",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"05"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"12",x"12",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"2d",x"2d",x"0d",x"0d",x"e8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"6d",x"51",x"4d",x"6d",x"51",x"4d",x"ac",x"c8",x"e8",x"c8",x"c8",x"c8",x"e8",x"e8",x"6d",x"89",x"c8",x"e8",x"e8",x"ec",x"ec",x"cc",x"4d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"29",x"2d",x"2e",x"32",x"32",x"32",x"32",x"32",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"2e",x"2d",x"09",x"09",x"09",x"09",x"25",x"24",x"09",x"09",x"09",x"09",x"2d",x"4d",x"49",x"49",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2d",x"2e",x"2e",x"2e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"29",x"91",x"90",x"6c",x"70",x"70",x"70",x"70",x"4d",x"2d",x"09",x"09",x"0a",x"0d",x"11",x"12",x"16",x"16",x"16",x"16",x"75",x"90",x"70",x"70",x"4c",x"4c",x"70",x"70",x"70",x"94",x"95",x"32",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2d",x"4d",x"6d",x"6d",x"6d",x"6d",x"29",x"49",x"6d",x"6d",x"4d",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"31",x"95",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"98",x"94",x"94",x"94",x"95",x"95",x"94",x"74",x"70",x"50",x"4c",x"50",x"71",x"50",x"4c",x"4c",x"50",x"50",x"51",x"50",x"50",x"51",x"4c",x"08",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0e",x"51",x"31",x"51",x"51",x"75",x"75",x"51",x"2d",x"51",x"51",x"51",x"51",x"50",x"50",x"70",x"90",x"70",x"6c",x"6c",x"70",x"6c",x"6c",x"90",x"91",x"94",x"98",x"98",x"95",x"4d",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"31",x"75",x"55",x"31",x"50",x"51",x"0d",x"09",x"09",x"09",x"8d",x"b5",x"91",x"6d",x"b1",x"95",x"30",x"55",x"75",x"75",x"51",x"50",x"75",x"31",x"0e",x"71",x"70",x"50",x"71",x"70",x"70",x"51",x"2d",x"2d",x"2d",x"2d",x"2c",x"2c",x"2c",x"08",x"08",x"04",x"2c",x"b8",x"fc",x"d8",x"70",x"b4",x"b4",x"4c",x"28",x"2c",x"2c",x"2c",x"50",x"74",x"75",x"75",x"74",x"70",x"2d",x"0d",x"05",x"05",x"09",x"09",x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"2d",x"8d",x"cc",x"ad",x"2d",x"0d",x"a8",x"c4",x"c4",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"a4",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"2d",x"49",x"a8",x"c8",x"c8",x"e8",x"e8",x"ec",x"ec",x"6d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"0d",x"0d",x"11",x"11",x"0d",x"29",x"29",x"2e",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4d",x"4d",x"4e",x"2e",x"32",x"32",x"52",x"2d",x"29",x"09",x"09",x"09",x"09",x"09",x"25",x"24",x"09",x"09",x"09",x"29",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"4d",x"4e",x"2e",x"2e",x"2e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"52",x"32",x"32",x"32",x"32",x"32",x"2e",x"29",x"94",x"70",x"70",x"70",x"70",x"71",x"70",x"09",x"09",x"09",x"0d",x"12",x"16",x"11",x"12",x"12",x"12",x"16",x"16",x"55",x"90",x"71",x"70",x"4c",x"4c",x"70",x"70",x"71",x"94",x"b4",x"75",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"4d",x"4d",x"4d",x"6d",x"4d",x"49",x"29",x"4d",x"6d",x"4d",x"2e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2d",x"71",x"98",x"b8",x"b9",x"b8",x"b8",x"b9",x"b8",x"b8",x"b8",x"98",x"98",x"98",x"98",x"94",x"94",x"95",x"95",x"95",x"94",x"94",x"75",x"71",x"4c",x"71",x"71",x"70",x"50",x"50",x"50",x"70",x"50",x"70",x"50",x"51",x"70",x"4d",x"28",x"28",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"2d",x"2d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"50",x"2c",x"2c",x"2c",x"70",x"90",x"70",x"6c",x"6c",x"70",x"6c",x"70",x"70",x"95",x"95",x"95",x"94",x"98",x"98",x"71",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"55",x"75",x"55",x"50",x"51",x"31",x"09",x"09",x"09",x"6d",x"b5",x"91",x"6d",x"91",x"b1",x"30",x"55",x"75",x"55",x"51",x"50",x"75",x"2d",x"2d",x"50",x"70",x"70",x"70",x"50",x"2d",x"31",x"31",x"2d",x"2d",x"2d",x"2d",x"2c",x"2c",x"08",x"08",x"08",x"08",x"4c",x"d8",x"fc",x"b4",x"70",x"b4",x"94",x"4c",x"2c",x"2c",x"2c",x"2d",x"50",x"50",x"50",x"50",x"2c",x"0d",x"09",x"09",x"05",x"09",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"09",x"05",x"09",x"09",x"11",x"12",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"4d",x"8d",x"ad",x"c8",x"e8",x"cc",x"4d",x"2d",x"ad",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"b1",x"88",x"a4",x"c4",x"c8",x"c8",x"c8",x"e8",x"ec",x"cc",x"6d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"16",x"11",x"11",x"0d",x"2d",x"2d",x"2d",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"32",x"32",x"32",x"32",x"52",x"4e",x"4d",x"4d",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"25",x"24",x"09",x"09",x"09",x"29",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"29",x"29",x"4d",x"4d",x"4d",x"4d",x"4d",x"2d",x"2d",x"2e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"29",x"6d",x"70",x"90",x"b4",x"94",x"70",x"70",x"51",x"0d",x"0d",x"11",x"12",x"12",x"16",x"15",x"12",x"12",x"12",x"12",x"16",x"36",x"90",x"70",x"70",x"4c",x"4c",x"4c",x"70",x"71",x"b4",x"b8",x"b9",x"75",x"55",x"36",x"16",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"4d",x"69",x"6d",x"4d",x"4d",x"49",x"29",x"49",x"6d",x"4d",x"2e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2d",x"71",x"94",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"99",x"99",x"98",x"94",x"95",x"95",x"94",x"95",x"95",x"74",x"70",x"71",x"71",x"75",x"75",x"74",x"51",x"51",x"70",x"70",x"70",x"70",x"50",x"51",x"50",x"51",x"2d",x"28",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"2e",x"2d",x"2d",x"51",x"51",x"51",x"2d",x"51",x"30",x"51",x"50",x"2c",x"2c",x"50",x"94",x"94",x"70",x"6c",x"6c",x"70",x"90",x"90",x"94",x"94",x"95",x"95",x"95",x"98",x"98",x"95",x"75",x"2d",x"0e",x"0e",x"0e",x"0e",x"0e",x"31",x"75",x"75",x"50",x"50",x"51",x"09",x"09",x"09",x"6d",x"b1",x"91",x"6d",x"8d",x"b1",x"51",x"55",x"75",x"75",x"51",x"51",x"75",x"31",x"4d",x"4c",x"71",x"70",x"74",x"71",x"0d",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2c",x"08",x"08",x"08",x"08",x"08",x"70",x"dc",x"dc",x"94",x"90",x"b4",x"70",x"2c",x"2c",x"2c",x"2d",x"2c",x"50",x"50",x"2d",x"0d",x"0d",x"09",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"05",x"09",x"0d",x"11",x"11",x"12",x"11",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"2d",x"6d",x"a8",x"e8",x"e8",x"e8",x"e8",x"cc",x"8d",x"8d",x"d0",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"c8",x"a4",x"a4",x"c4",x"c8",x"c8",x"c8",x"ec",x"ec",x"cc",x"4d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"15",x"11",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"0d",x"29",x"29",x"2d",x"2d",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2d",x"29",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"25",x"24",x"09",x"09",x"09",x"2d",x"4d",x"4d",x"2d",x"4d",x"4d",x"4d",x"4e",x"4d",x"4d",x"4d",x"4e",x"4e",x"4e",x"4e",x"2d",x"29",x"2d",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"2e",x"32",x"32",x"32",x"29",x"90",x"6c",x"94",x"d8",x"b4",x"94",x"70",x"51",x"12",x"12",x"16",x"16",x"12",x"12",x"12",x"11",x"12",x"12",x"12",x"12",x"35",x"b4",x"94",x"70",x"6c",x"4c",x"4c",x"70",x"95",x"b4",x"b4",x"b4",x"b4",x"b5",x"75",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4d",x"6d",x"6d",x"6d",x"4d",x"4d",x"29",x"29",x"4d",x"6d",x"4d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"12",x"12",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"51",x"94",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"98",x"98",x"98",x"94",x"94",x"94",x"94",x"94",x"75",x"70",x"70",x"75",x"75",x"75",x"71",x"70",x"50",x"71",x"70",x"70",x"51",x"50",x"51",x"50",x"50",x"51",x"2d",x"08",x"28",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0e",x"2d",x"2d",x"31",x"51",x"51",x"2d",x"51",x"30",x"51",x"51",x"50",x"50",x"90",x"d8",x"b4",x"90",x"6c",x"6c",x"70",x"94",x"b4",x"b4",x"b4",x"95",x"95",x"94",x"94",x"94",x"99",x"b8",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"75",x"79",x"54",x"50",x"51",x"2d",x"09",x"09",x"4d",x"91",x"b1",x"8d",x"6d",x"b1",x"71",x"55",x"75",x"75",x"51",x"51",x"75",x"51",x"4c",x"4c",x"71",x"74",x"95",x"51",x"09",x"09",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2c",x"08",x"08",x"08",x"28",x"05",x"08",x"94",x"dc",x"b8",x"90",x"94",x"94",x"4c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"0d",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"12",x"12",x"12",x"12",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"11",x"12",x"12",x"11",x"12",x"11",x"11",x"0d",x"11",x"11",x"11",x"11",x"11",x"0d",x"0d",x"89",x"e8",x"e8",x"e8",x"c8",x"c8",x"ec",x"ec",x"f0",x"f0",x"f0",x"c8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"cc",x"cc",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"c8",x"a4",x"a4",x"a4",x"c4",x"c4",x"c8",x"c8",x"e8",x"c8",x"8d",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"11",x"09",x"09",x"09",x"29",x"29",x"29",x"29",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"29",x"29",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"25",x"24",x"09",x"09",x"0d",x"2d",x"4d",x"4d",x"4d",x"4d",x"4d",x"2d",x"4e",x"4e",x"49",x"29",x"4e",x"4e",x"2e",x"2e",x"4e",x"4e",x"2d",x"29",x"2d",x"2e",x"2e",x"2e",x"32",x"2e",x"2e",x"2e",x"32",x"2e",x"32",x"32",x"2e",x"32",x"32",x"2d",x"6c",x"6c",x"94",x"b4",x"b8",x"b4",x"b4",x"94",x"71",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"55",x"b4",x"94",x"90",x"70",x"4c",x"4c",x"70",x"94",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"75",x"16",x"16",x"16",x"16",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"29",x"49",x"6d",x"6d",x"2e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"12",x"11",x"12",x"12",x"12",x"16",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"12",x"0e",x"0d",x"71",x"b8",x"b8",x"b8",x"98",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"98",x"98",x"94",x"94",x"94",x"94",x"71",x"70",x"70",x"75",x"95",x"74",x"74",x"74",x"71",x"50",x"70",x"70",x"70",x"71",x"51",x"71",x"50",x"50",x"4d",x"2d",x"09",x"28",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"2d",x"2d",x"31",x"2d",x"2d",x"51",x"51",x"51",x"51",x"51",x"71",x"b4",x"b4",x"b4",x"90",x"6c",x"6c",x"90",x"94",x"b4",x"b4",x"b4",x"b4",x"94",x"94",x"94",x"95",x"95",x"98",x"98",x"51",x"0e",x"0e",x"0e",x"0e",x"0e",x"75",x"79",x"75",x"51",x"51",x"31",x"09",x"09",x"4d",x"91",x"b1",x"8d",x"6d",x"b5",x"91",x"54",x"75",x"55",x"51",x"51",x"75",x"4d",x"4c",x"4c",x"70",x"94",x"71",x"0d",x"0d",x"09",x"09",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"08",x"09",x"09",x"09",x"09",x"08",x"28",x"b4",x"fc",x"94",x"71",x"94",x"94",x"2c",x"2c",x"2c",x"2c",x"2d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"0d",x"0d",x"0d",x"11",x"12",x"12",x"12",x"12",x"11",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"0d",x"0d",x"2d",x"89",x"e4",x"c4",x"c8",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"cc",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"a8",x"6d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"16",x"12",x"12",x"12",x"11",x"12",x"12",x"11",x"11",x"16",x"16",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"25",x"24",x"09",x"09",x"09",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"2d",x"2d",x"4d",x"49",x"29",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2e",x"2d",x"2d",x"2d",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"2d",x"4d",x"b4",x"70",x"b4",x"b8",x"b4",x"b4",x"b4",x"94",x"90",x"51",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"75",x"b8",x"b4",x"94",x"91",x"6c",x"4c",x"70",x"94",x"b4",x"b4",x"b4",x"b4",x"b8",x"b8",x"b5",x"36",x"16",x"1a",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"4d",x"8d",x"6d",x"4d",x"6d",x"6d",x"6d",x"49",x"29",x"49",x"6d",x"6d",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"12",x"12",x"0e",x"31",x"94",x"b8",x"b8",x"98",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"98",x"98",x"94",x"94",x"94",x"75",x"70",x"74",x"94",x"94",x"95",x"75",x"74",x"74",x"71",x"70",x"70",x"70",x"70",x"71",x"51",x"50",x"50",x"70",x"51",x"2d",x"09",x"28",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"2d",x"2d",x"2d",x"2d",x"4d",x"51",x"51",x"50",x"51",x"75",x"b5",x"b9",x"b4",x"b8",x"94",x"6c",x"6c",x"90",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"94",x"94",x"95",x"94",x"98",x"b8",x"75",x"31",x"0e",x"0e",x"0e",x"0e",x"51",x"99",x"79",x"51",x"51",x"55",x"0d",x"09",x"2d",x"91",x"b5",x"8d",x"6d",x"b1",x"91",x"55",x"55",x"55",x"51",x"50",x"75",x"4c",x"4c",x"6c",x"70",x"94",x"51",x"0e",x"0d",x"09",x"09",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"4d",x"b8",x"d8",x"94",x"90",x"b4",x"50",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"09",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"0d",x"0d",x"0d",x"69",x"e4",x"c8",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"ec",x"ec",x"f0",x"f0",x"f0",x"cc",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"88",x"2d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"11",x"15",x"11",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"24",x"25",x"09",x"09",x"09",x"49",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"2d",x"4d",x"4d",x"2d",x"2d",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"2e",x"2e",x"2d",x"2d",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2d",x"90",x"dc",x"70",x"b8",x"b8",x"b8",x"b8",x"b4",x"94",x"94",x"91",x"31",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"35",x"95",x"b8",x"b4",x"94",x"94",x"6c",x"4c",x"6c",x"94",x"b8",x"b4",x"94",x"b4",x"b8",x"b8",x"b8",x"75",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"8d",x"6d",x"4d",x"6d",x"6d",x"6d",x"4d",x"29",x"49",x"6d",x"6d",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"71",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"98",x"98",x"98",x"99",x"95",x"94",x"74",x"70",x"74",x"95",x"94",x"74",x"75",x"75",x"75",x"75",x"70",x"71",x"71",x"70",x"71",x"71",x"70",x"50",x"50",x"70",x"51",x"0d",x"09",x"28",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"31",x"51",x"2d",x"2d",x"4c",x"31",x"51",x"2c",x"51",x"95",x"d9",x"b9",x"b4",x"b8",x"94",x"6c",x"6c",x"90",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"94",x"95",x"94",x"98",x"99",x"98",x"51",x"0e",x"0e",x"0e",x"0e",x"2d",x"75",x"98",x"55",x"51",x"55",x"31",x"09",x"2d",x"91",x"b5",x"91",x"6d",x"91",x"b1",x"75",x"75",x"55",x"51",x"50",x"70",x"4c",x"4c",x"70",x"94",x"75",x"51",x"0e",x"09",x"09",x"09",x"09",x"0d",x"2d",x"2d",x"2d",x"09",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"71",x"d8",x"b4",x"70",x"94",x"95",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"0d",x"0d",x"11",x"12",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0e",x"4d",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"c8",x"c8",x"ec",x"e8",x"ec",x"f0",x"f0",x"f0",x"ec",x"cc",x"a8",x"a8",x"a4",x"a4",x"a8",x"c8",x"8d",x"2d",x"0e",x"0d",x"0d",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"12",x"16",x"11",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"24",x"29",x"0d",x"09",x"05",x"29",x"4d",x"4d",x"2d",x"4d",x"4d",x"4d",x"4d",x"4e",x"4d",x"4d",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"2e",x"32",x"32",x"2d",x"49",x"71",x"d8",x"d9",x"95",x"b5",x"d9",x"d9",x"d9",x"b4",x"90",x"94",x"90",x"70",x"51",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"55",x"b4",x"b4",x"b4",x"b4",x"94",x"70",x"4c",x"4c",x"94",x"b9",x"b8",x"b9",x"b8",x"b8",x"b8",x"b4",x"95",x"16",x"16",x"16",x"1a",x"16",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"6d",x"6d",x"6d",x"4d",x"6d",x"6d",x"49",x"29",x"49",x"6d",x"6d",x"2e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"71",x"b4",x"d8",x"b8",x"b8",x"98",x"b8",x"b8",x"98",x"98",x"99",x"95",x"95",x"74",x"94",x"95",x"94",x"95",x"74",x"74",x"75",x"75",x"75",x"70",x"70",x"70",x"71",x"71",x"70",x"51",x"51",x"50",x"94",x"71",x"09",x"09",x"28",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"28",x"31",x"51",x"51",x"51",x"2d",x"51",x"31",x"51",x"51",x"75",x"b9",x"d9",x"b9",x"b9",x"b8",x"94",x"6c",x"4c",x"90",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"94",x"94",x"99",x"98",x"98",x"98",x"71",x"2d",x"0e",x"0e",x"0e",x"0e",x"75",x"99",x"75",x"51",x"51",x"50",x"0d",x"09",x"91",x"b5",x"91",x"6d",x"91",x"b1",x"75",x"75",x"55",x"51",x"50",x"70",x"70",x"4c",x"71",x"90",x"71",x"2d",x"0e",x"09",x"0d",x"09",x"09",x"0d",x"0d",x"2d",x"09",x"08",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"b5",x"d8",x"94",x"70",x"b4",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"11",x"12",x"12",x"11",x"11",x"0d",x"0d",x"2d",x"4d",x"8d",x"ec",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"c8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"e8",x"e8",x"c8",x"ec",x"f0",x"f0",x"f0",x"ec",x"cc",x"cc",x"c8",x"c8",x"cc",x"ec",x"cc",x"8d",x"4d",x"0e",x"4d",x"89",x"6d",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"11",x"12",x"16",x"12",x"11",x"11",x"12",x"16",x"11",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"24",x"29",x"0d",x"09",x"24",x"29",x"2e",x"4e",x"4d",x"4d",x"4d",x"4d",x"4e",x"4e",x"4d",x"4d",x"4e",x"4e",x"2e",x"2e",x"4e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"2e",x"2d",x"2d",x"71",x"b4",x"d8",x"b9",x"95",x"90",x"b8",x"d9",x"b4",x"94",x"90",x"94",x"90",x"70",x"70",x"51",x"36",x"16",x"16",x"16",x"16",x"16",x"35",x"95",x"b4",x"b4",x"b4",x"b4",x"b4",x"90",x"4c",x"4c",x"70",x"b4",x"b8",x"b8",x"b8",x"b8",x"b5",x"94",x"75",x"16",x"16",x"16",x"1a",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"29",x"49",x"6d",x"6d",x"2e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"12",x"12",x"12",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"2d",x"71",x"94",x"b8",x"b8",x"b8",x"98",x"98",x"98",x"98",x"98",x"95",x"95",x"94",x"94",x"95",x"94",x"95",x"95",x"74",x"74",x"75",x"74",x"75",x"71",x"70",x"70",x"71",x"50",x"51",x"71",x"94",x"94",x"4d",x"0e",x"09",x"28",x"09",x"09",x"09",x"09",x"0d",x"0d",x"2d",x"2c",x"4c",x"51",x"51",x"51",x"51",x"51",x"31",x"51",x"51",x"95",x"d9",x"b9",x"b9",x"b9",x"b9",x"b5",x"6c",x"4c",x"90",x"b4",x"b8",x"b4",x"b4",x"b8",x"d8",x"b8",x"95",x"94",x"98",x"99",x"98",x"99",x"75",x"2d",x"0e",x"0e",x"0e",x"0a",x"51",x"99",x"75",x"51",x"30",x"54",x"31",x"09",x"6d",x"b5",x"91",x"6d",x"91",x"b1",x"95",x"75",x"55",x"50",x"50",x"70",x"50",x"4c",x"71",x"94",x"71",x"2d",x"0e",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"4d",x"b8",x"d8",x"90",x"94",x"71",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"0d",x"12",x"12",x"12",x"11",x"11",x"0d",x"0d",x"6d",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"ec",x"c8",x"ec",x"c8",x"a4",x"a4",x"a4",x"a8",x"a4",x"a8",x"84",x"a4",x"a8",x"c8",x"e8",x"c8",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ad",x"2d",x"89",x"e4",x"e8",x"ad",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"12",x"16",x"16",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"24",x"09",x"0d",x"0d",x"24",x"25",x"31",x"32",x"4e",x"4d",x"4d",x"4d",x"4e",x"4e",x"4d",x"4d",x"4d",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"29",x"29",x"2d",x"95",x"d8",x"b4",x"b4",x"94",x"6c",x"94",x"b4",x"94",x"90",x"94",x"94",x"71",x"70",x"70",x"70",x"55",x"16",x"16",x"16",x"16",x"16",x"55",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"95",x"6c",x"4c",x"6c",x"94",x"b9",x"b4",x"b8",x"b4",x"95",x"94",x"55",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"2e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"09",x"09",x"0d",x"11",x"16",x"16",x"16",x"16",x"16",x"12",x"11",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"12",x"12",x"0e",x"0d",x"51",x"94",x"b8",x"b8",x"98",x"98",x"99",x"98",x"98",x"98",x"95",x"95",x"95",x"95",x"95",x"95",x"95",x"94",x"74",x"74",x"74",x"75",x"71",x"70",x"70",x"70",x"50",x"71",x"94",x"94",x"4c",x"09",x"0e",x"0d",x"28",x"08",x"09",x"09",x"09",x"0d",x"2d",x"4c",x"4c",x"4c",x"51",x"51",x"51",x"51",x"51",x"51",x"2c",x"31",x"95",x"d9",x"b9",x"b9",x"b9",x"b9",x"b9",x"71",x"4c",x"90",x"b4",x"b8",x"b8",x"b8",x"b9",x"d9",x"b9",x"99",x"98",x"98",x"99",x"98",x"98",x"74",x"2d",x"0e",x"0e",x"0e",x"0e",x"31",x"75",x"79",x"54",x"30",x"55",x"75",x"09",x"6d",x"b1",x"91",x"6d",x"6d",x"91",x"91",x"75",x"55",x"50",x"50",x"70",x"50",x"51",x"50",x"70",x"51",x"2d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"75",x"fc",x"b4",x"70",x"b4",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"05",x"09",x"11",x"11",x"11",x"12",x"11",x"0e",x"31",x"ad",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"f0",x"f0",x"c8",x"e8",x"c8",x"a4",x"84",x"88",x"84",x"a4",x"88",x"88",x"84",x"a8",x"c8",x"ec",x"ec",x"cc",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"ec",x"cc",x"c8",x"c8",x"ec",x"ec",x"ec",x"ac",x"a8",x"c4",x"e4",x"e8",x"a8",x"4d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"16",x"16",x"12",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"24",x"09",x"0d",x"0d",x"24",x"29",x"09",x"2d",x"52",x"52",x"4e",x"4d",x"4d",x"4d",x"4e",x"4e",x"2e",x"4e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"2d",x"29",x"2d",x"0d",x"12",x"51",x"95",x"b4",x"94",x"94",x"6c",x"6c",x"71",x"94",x"90",x"90",x"71",x"71",x"70",x"70",x"71",x"36",x"16",x"16",x"16",x"12",x"12",x"75",x"b8",x"b4",x"b4",x"b4",x"94",x"b8",x"95",x"70",x"4c",x"4c",x"95",x"95",x"b4",x"95",x"95",x"90",x"70",x"55",x"16",x"16",x"16",x"16",x"16",x"16",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"6d",x"91",x"91",x"6d",x"69",x"6d",x"6d",x"4d",x"29",x"29",x"6d",x"6d",x"2e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"12",x"12",x"11",x"11",x"11",x"12",x"11",x"11",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"4d",x"70",x"94",x"b8",x"b8",x"b8",x"b8",x"94",x"94",x"94",x"94",x"94",x"95",x"95",x"95",x"95",x"94",x"74",x"74",x"75",x"71",x"71",x"51",x"51",x"74",x"95",x"b4",x"90",x"4d",x"09",x"0d",x"0e",x"0d",x"08",x"08",x"09",x"09",x"09",x"0d",x"4d",x"50",x"50",x"4c",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"30",x"95",x"d9",x"d9",x"b9",x"d9",x"dd",x"b9",x"71",x"6d",x"91",x"b5",x"b9",x"b9",x"b9",x"b5",x"95",x"95",x"98",x"99",x"98",x"99",x"98",x"98",x"71",x"2d",x"0e",x"0e",x"0e",x"0e",x"0d",x"55",x"78",x"55",x"31",x"55",x"75",x"0d",x"6d",x"91",x"91",x"6d",x"6d",x"91",x"91",x"55",x"55",x"51",x"51",x"50",x"51",x"51",x"30",x"30",x"30",x"30",x"51",x"75",x"2d",x"09",x"0a",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"2d",x"94",x"fc",x"90",x"94",x"51",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"0d",x"12",x"12",x"12",x"12",x"12",x"4d",x"91",x"ec",x"ec",x"e8",x"c8",x"c8",x"c8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"c8",x"c8",x"c8",x"a4",x"84",x"84",x"84",x"84",x"84",x"84",x"a8",x"c8",x"ec",x"ec",x"c8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a8",x"a8",x"c8",x"c8",x"e8",x"ec",x"c8",x"c4",x"c4",x"e8",x"e8",x"ad",x"4d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"16",x"16",x"12",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"04",x"24",x"09",x"0d",x"0d",x"24",x"29",x"09",x"0d",x"2d",x"2e",x"52",x"2e",x"2e",x"4e",x"4e",x"2e",x"4e",x"4e",x"2e",x"2e",x"2e",x"4e",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2d",x"2d",x"2c",x"31",x"12",x"12",x"11",x"51",x"75",x"94",x"94",x"70",x"4c",x"70",x"90",x"90",x"70",x"70",x"70",x"70",x"70",x"51",x"16",x"16",x"12",x"12",x"12",x"12",x"75",x"b8",x"b5",x"94",x"b4",x"b4",x"b9",x"95",x"70",x"4c",x"4c",x"70",x"94",x"94",x"95",x"71",x"70",x"70",x"36",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"2e",x"4d",x"91",x"95",x"91",x"6d",x"6d",x"6d",x"49",x"29",x"29",x"6d",x"6d",x"4d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"12",x"12",x"12",x"16",x"16",x"12",x"16",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"2d",x"51",x"94",x"b4",x"b8",x"b8",x"b8",x"b8",x"98",x"94",x"95",x"94",x"94",x"95",x"75",x"75",x"74",x"75",x"75",x"74",x"94",x"95",x"95",x"94",x"94",x"90",x"4c",x"09",x"09",x"0d",x"0d",x"0d",x"08",x"08",x"09",x"09",x"09",x"2d",x"50",x"50",x"50",x"50",x"50",x"51",x"51",x"51",x"51",x"71",x"51",x"50",x"95",x"d9",x"d9",x"d9",x"d9",x"dd",x"b9",x"71",x"71",x"71",x"b5",x"b9",x"b5",x"95",x"95",x"95",x"95",x"98",x"98",x"99",x"98",x"98",x"74",x"51",x"0d",x"0e",x"0d",x"0e",x"0e",x"09",x"55",x"78",x"75",x"31",x"51",x"75",x"31",x"6d",x"91",x"91",x"8d",x"6d",x"91",x"91",x"75",x"55",x"51",x"51",x"31",x"51",x"51",x"51",x"30",x"30",x"50",x"50",x"75",x"71",x"51",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"51",x"d8",x"d8",x"90",x"95",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"0d",x"11",x"12",x"12",x"12",x"32",x"b1",x"ec",x"ec",x"c8",x"c8",x"c8",x"a8",x"a8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"c8",x"c8",x"c8",x"a4",x"84",x"84",x"a4",x"84",x"84",x"a8",x"c8",x"ec",x"ec",x"c8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"ec",x"c8",x"a8",x"84",x"a8",x"a8",x"c8",x"e8",x"cc",x"c8",x"c8",x"c8",x"e8",x"e8",x"ac",x"0d",x"0d",x"0d",x"0d",x"11",x"16",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"16",x"16",x"12",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"24",x"24",x"09",x"0d",x"0d",x"24",x"29",x"0d",x"09",x"29",x"29",x"2e",x"32",x"32",x"32",x"32",x"2e",x"4e",x"4e",x"2e",x"2e",x"4e",x"4e",x"2e",x"2e",x"52",x"32",x"32",x"32",x"32",x"29",x"29",x"29",x"50",x"54",x"31",x"12",x"11",x"11",x"11",x"31",x"71",x"90",x"95",x"70",x"6c",x"70",x"71",x"71",x"70",x"70",x"70",x"71",x"31",x"12",x"12",x"12",x"12",x"12",x"32",x"75",x"b8",x"94",x"94",x"b5",x"b8",x"b8",x"95",x"94",x"70",x"48",x"4c",x"70",x"70",x"70",x"70",x"70",x"75",x"16",x"16",x"16",x"16",x"12",x"11",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"2e",x"4d",x"6d",x"91",x"91",x"91",x"6d",x"6d",x"4d",x"29",x"49",x"6d",x"6d",x"4d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"11",x"0d",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"0e",x"0d",x"2d",x"50",x"94",x"b8",x"b8",x"b8",x"b8",x"98",x"95",x"94",x"94",x"95",x"95",x"95",x"95",x"75",x"74",x"94",x"b4",x"b8",x"b8",x"94",x"70",x"2c",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"28",x"08",x"09",x"09",x"09",x"2d",x"50",x"50",x"51",x"50",x"50",x"71",x"75",x"51",x"51",x"75",x"75",x"75",x"95",x"b9",x"d9",x"d9",x"d9",x"d9",x"b9",x"95",x"71",x"71",x"95",x"95",x"95",x"95",x"95",x"95",x"99",x"98",x"98",x"99",x"98",x"98",x"74",x"2d",x"0d",x"0e",x"09",x"0e",x"0e",x"09",x"31",x"79",x"75",x"51",x"31",x"55",x"55",x"71",x"91",x"91",x"6d",x"6d",x"91",x"91",x"75",x"55",x"55",x"51",x"51",x"2c",x"51",x"51",x"55",x"51",x"51",x"51",x"30",x"75",x"99",x"51",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"75",x"fc",x"94",x"b4",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"12",x"71",x"ac",x"ad",x"71",x"b1",x"ec",x"ec",x"e8",x"c8",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"e8",x"c8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"c4",x"c8",x"c8",x"c8",x"a8",x"a8",x"c8",x"c8",x"c8",x"ec",x"ec",x"c8",x"a8",x"a8",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"c8",x"c8",x"a8",x"84",x"a8",x"a4",x"a8",x"c8",x"ec",x"cc",x"c8",x"c8",x"c8",x"e8",x"e8",x"8d",x"11",x"11",x"0d",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"16",x"16",x"11",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"24",x"25",x"09",x"0d",x"0d",x"24",x"29",x"0d",x"09",x"09",x"09",x"29",x"29",x"2d",x"2d",x"4e",x"52",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"29",x"29",x"29",x"29",x"2d",x"31",x"31",x"51",x"50",x"11",x"12",x"12",x"12",x"12",x"12",x"31",x"71",x"70",x"70",x"4c",x"4c",x"71",x"71",x"70",x"70",x"70",x"31",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"75",x"d8",x"b8",x"b8",x"b9",x"b8",x"b8",x"94",x"71",x"70",x"48",x"4c",x"70",x"71",x"70",x"70",x"71",x"51",x"16",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0e",x"0e",x"0d",x"4d",x"4d",x"6d",x"91",x"91",x"91",x"91",x"6d",x"29",x"4d",x"6d",x"6d",x"4d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"31",x"51",x"70",x"70",x"94",x"b4",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b8",x"b4",x"b8",x"94",x"94",x"70",x"6c",x"4d",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"28",x"08",x"09",x"09",x"09",x"2d",x"50",x"50",x"50",x"51",x"50",x"50",x"71",x"71",x"51",x"75",x"75",x"75",x"75",x"95",x"b9",x"b5",x"b5",x"99",x"95",x"75",x"71",x"71",x"71",x"75",x"95",x"95",x"95",x"95",x"98",x"99",x"98",x"98",x"99",x"b8",x"51",x"0d",x"09",x"0d",x"09",x"0d",x"0e",x"09",x"2d",x"75",x"79",x"55",x"30",x"55",x"75",x"71",x"91",x"91",x"6d",x"49",x"91",x"91",x"75",x"55",x"51",x"31",x"30",x"55",x"75",x"75",x"79",x"75",x"55",x"55",x"55",x"54",x"75",x"99",x"51",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"2d",x"b8",x"d8",x"b4",x"51",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"71",x"cd",x"e8",x"ec",x"cc",x"ec",x"ec",x"ec",x"c8",x"a8",x"a8",x"a8",x"a8",x"a4",x"a8",x"c8",x"c8",x"a8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"c4",x"c8",x"e8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"c8",x"c8",x"a8",x"a8",x"ec",x"ec",x"ec",x"ec",x"cc",x"c8",x"e8",x"c8",x"a8",x"84",x"84",x"84",x"84",x"a8",x"cc",x"cc",x"cc",x"c8",x"c8",x"e8",x"e8",x"ad",x"11",x"12",x"11",x"11",x"12",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"16",x"12",x"11",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"24",x"25",x"09",x"0d",x"0d",x"24",x"29",x"0d",x"09",x"09",x"09",x"09",x"09",x"29",x"29",x"2d",x"2d",x"2d",x"2d",x"2e",x"2e",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"29",x"2d",x"2c",x"50",x"50",x"51",x"51",x"51",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"31",x"71",x"70",x"4c",x"4c",x"4c",x"71",x"70",x"70",x"70",x"31",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"55",x"b9",x"b8",x"b8",x"b9",x"b8",x"94",x"90",x"70",x"70",x"4c",x"4c",x"4c",x"71",x"70",x"70",x"71",x"51",x"0e",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0d",x"49",x"49",x"49",x"6d",x"91",x"91",x"91",x"6d",x"4d",x"71",x"8d",x"6d",x"4d",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"2d",x"31",x"51",x"71",x"70",x"90",x"94",x"94",x"94",x"94",x"90",x"90",x"94",x"70",x"4d",x"2d",x"2d",x"09",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0d",x"28",x"09",x"09",x"09",x"09",x"2d",x"50",x"50",x"50",x"51",x"51",x"50",x"70",x"51",x"51",x"51",x"75",x"75",x"75",x"75",x"95",x"95",x"95",x"95",x"95",x"71",x"71",x"4d",x"71",x"71",x"95",x"95",x"95",x"98",x"98",x"99",x"99",x"98",x"b8",x"94",x"2d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"0d",x"55",x"79",x"55",x"31",x"51",x"55",x"75",x"91",x"91",x"6d",x"49",x"91",x"91",x"75",x"55",x"31",x"30",x"51",x"75",x"79",x"79",x"79",x"75",x"75",x"55",x"75",x"55",x"55",x"78",x"75",x"51",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"71",x"d8",x"b4",x"95",x"2d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"cc",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"c8",x"a8",x"a8",x"a4",x"a4",x"88",x"84",x"c8",x"e8",x"c8",x"a8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"a8",x"a4",x"c4",x"c8",x"e8",x"c8",x"c8",x"e8",x"e8",x"e8",x"c8",x"c8",x"a4",x"a8",x"cc",x"ec",x"ec",x"ec",x"ec",x"c8",x"c4",x"e8",x"c8",x"a8",x"a4",x"84",x"a4",x"84",x"84",x"c8",x"e8",x"cc",x"c8",x"c8",x"e8",x"e8",x"91",x"12",x"12",x"11",x"12",x"12",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"12",x"11",x"12",x"16",x"12",x"11",x"0d",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"24",x"05",x"09",x"0d",x"0d",x"24",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"29",x"09",x"29",x"29",x"29",x"29",x"2d",x"50",x"50",x"50",x"55",x"51",x"51",x"51",x"50",x"50",x"50",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"51",x"70",x"70",x"4c",x"4c",x"70",x"71",x"70",x"90",x"31",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"75",x"b4",x"b4",x"94",x"94",x"71",x"70",x"70",x"70",x"4c",x"4c",x"4c",x"50",x"50",x"70",x"70",x"51",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"2d",x"49",x"4d",x"4d",x"49",x"6d",x"6d",x"6d",x"6d",x"71",x"b5",x"91",x"6d",x"4d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"29",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"28",x"09",x"09",x"09",x"09",x"2c",x"50",x"51",x"51",x"50",x"50",x"70",x"70",x"50",x"51",x"51",x"75",x"75",x"75",x"75",x"74",x"75",x"95",x"95",x"75",x"71",x"71",x"71",x"71",x"71",x"71",x"95",x"95",x"98",x"98",x"99",x"99",x"b8",x"94",x"4d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"51",x"78",x"54",x"31",x"31",x"55",x"75",x"91",x"91",x"8d",x"49",x"91",x"95",x"75",x"51",x"2d",x"30",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"31",x"75",x"55",x"31",x"55",x"99",x"74",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"95",x"b8",x"b4",x"31",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"88",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"cc",x"c8",x"a8",x"a8",x"84",x"84",x"84",x"a4",x"c8",x"c8",x"c8",x"a8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"a8",x"a4",x"a4",x"c4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"a4",x"a8",x"cc",x"ec",x"ec",x"ec",x"cc",x"c8",x"a4",x"c8",x"c8",x"c8",x"a8",x"a8",x"84",x"84",x"84",x"a8",x"e8",x"c8",x"c8",x"c8",x"c8",x"8d",x"11",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"16",x"16",x"16",x"11",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"24",x"05",x"09",x"09",x"0d",x"25",x"25",x"09",x"0d",x"09",x"09",x"09",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"11",x"51",x"50",x"50",x"51",x"51",x"55",x"55",x"55",x"75",x"51",x"31",x"31",x"50",x"50",x"50",x"11",x"12",x"11",x"11",x"12",x"11",x"12",x"12",x"11",x"71",x"90",x"70",x"4c",x"70",x"91",x"70",x"90",x"51",x"12",x"12",x"12",x"12",x"12",x"31",x"11",x"12",x"12",x"55",x"75",x"71",x"90",x"90",x"70",x"70",x"71",x"4c",x"48",x"4c",x"50",x"70",x"70",x"70",x"70",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0d",x"2d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"29",x"29",x"6d",x"6d",x"6d",x"6d",x"2e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"28",x"08",x"09",x"09",x"09",x"2c",x"51",x"50",x"50",x"50",x"51",x"50",x"50",x"70",x"71",x"51",x"75",x"75",x"75",x"75",x"75",x"75",x"95",x"95",x"71",x"71",x"71",x"71",x"71",x"71",x"71",x"95",x"95",x"99",x"98",x"b8",x"b8",x"94",x"51",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"31",x"79",x"75",x"51",x"31",x"55",x"55",x"71",x"91",x"91",x"49",x"91",x"75",x"55",x"31",x"30",x"51",x"75",x"75",x"75",x"74",x"74",x"74",x"51",x"2d",x"0d",x"2d",x"31",x"51",x"75",x"98",x"75",x"31",x"0e",x"11",x"0e",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"32",x"d8",x"b4",x"75",x"31",x"0d",x"0d",x"0d",x"11",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"11",x"0d",x"0d",x"0d",x"11",x"11"),
(x"09",x"05",x"05",x"09",x"05",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"05",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"c8",x"e8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"a8",x"a8",x"84",x"84",x"88",x"a8",x"c8",x"e8",x"c8",x"c8",x"a8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"c8",x"a8",x"a4",x"a4",x"a4",x"c4",x"c4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"c8",x"cc",x"ec",x"ec",x"ec",x"cc",x"a8",x"a4",x"c4",x"c8",x"c8",x"c8",x"a8",x"a8",x"a4",x"a4",x"c8",x"e8",x"c8",x"c8",x"c8",x"a8",x"6d",x"11",x"12",x"11",x"11",x"12",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"11",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"29",x"29",x"29",x"09",x"29",x"25",x"09",x"09",x"09",x"0d",x"25",x"24",x"09",x"0d",x"09",x"09",x"29",x"4d",x"4e",x"4d",x"4e",x"4e",x"2e",x"2e",x"32",x"55",x"55",x"54",x"54",x"55",x"75",x"75",x"75",x"55",x"50",x"30",x"31",x"51",x"51",x"50",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"12",x"12",x"51",x"95",x"70",x"6c",x"70",x"95",x"94",x"94",x"95",x"51",x"31",x"31",x"31",x"31",x"51",x"51",x"31",x"11",x"12",x"35",x"55",x"51",x"71",x"90",x"70",x"70",x"50",x"4c",x"48",x"4c",x"70",x"70",x"70",x"94",x"51",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"2d",x"4d",x"4d",x"49",x"4d",x"4d",x"49",x"25",x"05",x"29",x"6d",x"4d",x"49",x"4d",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"28",x"09",x"09",x"09",x"09",x"4c",x"71",x"50",x"50",x"50",x"51",x"50",x"51",x"70",x"70",x"51",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"95",x"71",x"71",x"71",x"71",x"71",x"71",x"71",x"95",x"95",x"99",x"98",x"94",x"94",x"51",x"0d",x"0e",x"12",x"12",x"12",x"11",x"12",x"12",x"12",x"11",x"0e",x"31",x"75",x"75",x"51",x"30",x"51",x"55",x"75",x"91",x"8d",x"49",x"91",x"75",x"55",x"30",x"30",x"55",x"75",x"75",x"74",x"70",x"70",x"55",x"51",x"2d",x"09",x"0d",x"2d",x"31",x"51",x"98",x"99",x"51",x"12",x"12",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"31",x"31",x"31",x"31",x"31",x"31",x"b8",x"d8",x"b4",x"51",x"0d",x"0d",x"0d",x"0d",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"0d",x"0d",x"0d",x"11",x"12"),
(x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"69",x"e8",x"c8",x"ec",x"ec",x"ec",x"ec",x"e8",x"ec",x"c8",x"a4",x"84",x"84",x"a8",x"c8",x"e8",x"c8",x"c8",x"a4",x"a8",x"c8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"c8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"c8",x"cc",x"ec",x"ec",x"ec",x"ec",x"cc",x"a8",x"a4",x"a4",x"c4",x"c4",x"c8",x"e8",x"e8",x"c8",x"c8",x"e8",x"e8",x"c8",x"c8",x"ac",x"c8",x"c8",x"71",x"12",x"51",x"71",x"51",x"12",x"16",x"12",x"11",x"11",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"2e",x"2e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4d",x"29",x"09",x"09",x"09",x"0d",x"29",x"24",x"09",x"09",x"09",x"09",x"49",x"49",x"29",x"29",x"4d",x"4d",x"2d",x"2e",x"2e",x"2e",x"31",x"55",x"54",x"51",x"75",x"55",x"55",x"55",x"51",x"31",x"31",x"51",x"51",x"50",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"12",x"12",x"31",x"75",x"90",x"6c",x"70",x"b4",x"b8",x"b8",x"b4",x"94",x"90",x"90",x"70",x"6c",x"70",x"70",x"70",x"71",x"35",x"16",x"16",x"16",x"55",x"91",x"70",x"70",x"70",x"4c",x"48",x"4c",x"4c",x"70",x"70",x"94",x"b5",x"51",x"0d",x"09",x"09",x"0d",x"0d",x"0e",x"0d",x"2e",x"4d",x"4d",x"4d",x"4d",x"49",x"4d",x"49",x"05",x"05",x"29",x"4d",x"4d",x"6d",x"6d",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"28",x"09",x"09",x"09",x"09",x"4c",x"94",x"70",x"50",x"4c",x"50",x"51",x"51",x"50",x"50",x"71",x"71",x"74",x"75",x"75",x"75",x"75",x"75",x"95",x"75",x"71",x"71",x"71",x"51",x"71",x"71",x"95",x"b9",x"b9",x"b9",x"74",x"2d",x"0d",x"0d",x"12",x"12",x"0e",x"0d",x"12",x"11",x"11",x"0d",x"11",x"0e",x"31",x"75",x"75",x"55",x"30",x"31",x"55",x"75",x"91",x"8d",x"49",x"71",x"55",x"55",x"31",x"51",x"75",x"75",x"75",x"70",x"90",x"71",x"51",x"71",x"51",x"0e",x"0d",x"09",x"08",x"2d",x"75",x"b8",x"95",x"31",x"0e",x"12",x"0d",x"31",x"31",x"31",x"51",x"51",x"51",x"74",x"75",x"75",x"75",x"55",x"75",x"95",x"d8",x"b4",x"51",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"12",x"0d",x"0d",x"11",x"11",x"12"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"45",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"ec",x"c8",x"c8",x"a8",x"c8",x"c8",x"e8",x"e8",x"c8",x"c8",x"a4",x"a8",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a4",x"a8",x"a8",x"a8",x"a8",x"c8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"a8",x"a4",x"a4",x"a4",x"c4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"cc",x"a8",x"c8",x"c8",x"ac",x"8d",x"ac",x"cc",x"cc",x"ad",x"4d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"2e",x"2e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4d",x"29",x"09",x"09",x"09",x"0d",x"29",x"24",x"09",x"09",x"09",x"09",x"49",x"29",x"29",x"29",x"29",x"29",x"2e",x"2e",x"2e",x"2e",x"32",x"31",x"51",x"55",x"54",x"55",x"55",x"55",x"51",x"31",x"31",x"31",x"51",x"50",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"32",x"75",x"94",x"90",x"4c",x"b8",x"b4",x"b8",x"b8",x"94",x"90",x"90",x"70",x"70",x"70",x"70",x"70",x"70",x"51",x"16",x"16",x"1a",x"16",x"51",x"70",x"50",x"70",x"6c",x"4c",x"4c",x"4c",x"50",x"74",x"98",x"b8",x"94",x"71",x"51",x"0d",x"09",x"0d",x"0d",x"2d",x"49",x"6d",x"4d",x"4d",x"4d",x"4d",x"49",x"05",x"05",x"29",x"49",x"4d",x"4d",x"4d",x"2e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"16",x"16",x"16",x"12",x"12",x"12",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"28",x"09",x"09",x"09",x"08",x"28",x"51",x"94",x"95",x"50",x"51",x"51",x"50",x"50",x"71",x"70",x"71",x"74",x"75",x"75",x"75",x"75",x"75",x"74",x"95",x"75",x"71",x"71",x"4d",x"71",x"71",x"95",x"b9",x"b9",x"b9",x"95",x"51",x"0a",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"11",x"51",x"74",x"55",x"2c",x"31",x"55",x"55",x"71",x"8d",x"69",x"75",x"55",x"31",x"31",x"51",x"75",x"75",x"70",x"70",x"90",x"71",x"51",x"51",x"51",x"31",x"0e",x"08",x"08",x"08",x"50",x"98",x"b9",x"51",x"31",x"31",x"31",x"31",x"31",x"4d",x"51",x"51",x"51",x"50",x"51",x"51",x"30",x"31",x"75",x"75",x"95",x"b4",x"71",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"12",x"11",x"11",x"12",x"16",x"12"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"05",x"09",x"09",x"09",x"05",x"09",x"09",x"05",x"09",x"09",x"09",x"25",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"c8",x"c8",x"a4",x"a4",x"c8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"cc",x"c8",x"a8",x"a8",x"a8",x"a8",x"c8",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c8",x"a4",x"c8",x"cc",x"cc",x"a8",x"c8",x"c8",x"c8",x"e8",x"ec",x"e8",x"e8",x"e8",x"a8",x"29",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0d",x"2e",x"4e",x"4e",x"4e",x"4e",x"4e",x"2d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"29",x"09",x"09",x"0d",x"09",x"24",x"09",x"09",x"09",x"09",x"25",x"29",x"29",x"29",x"29",x"29",x"2e",x"2e",x"2e",x"32",x"32",x"2e",x"31",x"51",x"54",x"55",x"55",x"55",x"51",x"31",x"31",x"31",x"51",x"50",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"75",x"b8",x"94",x"4c",x"94",x"b4",x"b9",x"b8",x"94",x"74",x"74",x"70",x"70",x"70",x"70",x"70",x"70",x"70",x"35",x"16",x"16",x"12",x"31",x"70",x"70",x"50",x"70",x"4c",x"48",x"4c",x"70",x"74",x"94",x"94",x"b8",x"b8",x"95",x"51",x"0d",x"0d",x"0d",x"4d",x"69",x"69",x"4d",x"4d",x"4d",x"4d",x"25",x"05",x"29",x"4d",x"4d",x"4d",x"4d",x"2d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"28",x"09",x"09",x"09",x"08",x"08",x"0d",x"70",x"94",x"74",x"71",x"71",x"50",x"50",x"71",x"70",x"70",x"70",x"75",x"75",x"75",x"75",x"75",x"75",x"95",x"95",x"75",x"71",x"4d",x"71",x"95",x"95",x"b9",x"b9",x"b9",x"b9",x"75",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"11",x"0d",x"31",x"75",x"75",x"30",x"31",x"55",x"55",x"75",x"8d",x"6d",x"55",x"55",x"31",x"51",x"55",x"75",x"75",x"6c",x"71",x"70",x"71",x"51",x"50",x"51",x"51",x"0d",x"08",x"04",x"08",x"2c",x"95",x"d9",x"75",x"71",x"2d",x"2c",x"2c",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"0c",x"31",x"74",x"75",x"36",x"95",x"95",x"11",x"0e",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"0d"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"29",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"a4",x"a4",x"a8",x"c8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"cc",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"c8",x"ec",x"cc",x"a8",x"c8",x"c8",x"c8",x"ec",x"ec",x"c8",x"a8",x"c8",x"e8",x"c8",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"2e",x"32",x"2e",x"2e",x"4e",x"4e",x"4e",x"4e",x"4d",x"29",x"29",x"29",x"29",x"29",x"49",x"29",x"09",x"09",x"09",x"0d",x"24",x"09",x"09",x"09",x"09",x"25",x"29",x"29",x"29",x"29",x"29",x"29",x"2e",x"2e",x"2e",x"32",x"32",x"2e",x"31",x"54",x"55",x"55",x"55",x"51",x"31",x"31",x"31",x"30",x"50",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"11",x"12",x"75",x"b8",x"94",x"4c",x"90",x"b9",x"b9",x"b8",x"94",x"94",x"74",x"70",x"70",x"70",x"70",x"70",x"70",x"70",x"51",x"16",x"11",x"09",x"2d",x"71",x"70",x"51",x"50",x"4c",x"48",x"4c",x"70",x"94",x"94",x"95",x"95",x"98",x"b8",x"b5",x"51",x"0d",x"31",x"49",x"69",x"49",x"4d",x"6d",x"4d",x"29",x"05",x"29",x"4d",x"4d",x"4d",x"4d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"28",x"09",x"09",x"09",x"08",x"08",x"0d",x"09",x"70",x"94",x"94",x"94",x"70",x"51",x"50",x"51",x"70",x"51",x"71",x"75",x"75",x"74",x"75",x"99",x"b9",x"95",x"95",x"71",x"4d",x"51",x"95",x"b9",x"b9",x"b9",x"b5",x"b9",x"b9",x"75",x"09",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"0d",x"0d",x"11",x"0d",x"0e",x"31",x"75",x"55",x"31",x"31",x"51",x"55",x"75",x"8d",x"6d",x"55",x"55",x"31",x"51",x"55",x"75",x"75",x"6c",x"71",x"70",x"51",x"51",x"50",x"50",x"50",x"0d",x"04",x"08",x"08",x"0d",x"75",x"dc",x"74",x"95",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"0d",x"0d",x"50",x"74",x"74",x"31",x"12",x"55",x"95",x"51",x"0e",x"12",x"12",x"0d",x"12",x"12",x"12",x"11",x"12",x"12",x"12",x"11",x"0d",x"0d",x"09",x"05",x"05"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"0d",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"49",x"88",x"ac",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"c8",x"c8",x"c4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"a8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"cc",x"ec",x"cc",x"a8",x"a8",x"a8",x"c8",x"ec",x"ec",x"c8",x"a4",x"a8",x"c8",x"e8",x"a8",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"2e",x"32",x"52",x"4e",x"2e",x"2e",x"4e",x"4d",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"09",x"09",x"09",x"0d",x"24",x"09",x"09",x"09",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2e",x"2e",x"2e",x"32",x"32",x"32",x"2e",x"2d",x"54",x"55",x"55",x"55",x"51",x"31",x"31",x"31",x"30",x"50",x"11",x"11",x"11",x"12",x"12",x"11",x"12",x"12",x"11",x"12",x"75",x"b8",x"94",x"70",x"70",x"b9",x"b8",x"94",x"70",x"70",x"70",x"50",x"70",x"70",x"70",x"70",x"70",x"70",x"71",x"0d",x"0d",x"09",x"2d",x"71",x"70",x"70",x"70",x"71",x"4c",x"48",x"4c",x"74",x"94",x"94",x"94",x"94",x"98",x"b8",x"75",x"2d",x"51",x"49",x"4d",x"49",x"49",x"6d",x"49",x"05",x"05",x"4d",x"4d",x"49",x"4d",x"2d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"29",x"28",x"09",x"09",x"09",x"28",x"28",x"0e",x"09",x"2d",x"4c",x"70",x"90",x"94",x"94",x"94",x"94",x"95",x"95",x"74",x"94",x"95",x"94",x"95",x"99",x"b9",x"b9",x"95",x"95",x"51",x"4d",x"75",x"b9",x"b9",x"b9",x"b9",x"b9",x"d9",x"b9",x"0d",x"0d",x"09",x"0d",x"09",x"09",x"0e",x"12",x"12",x"11",x"12",x"12",x"11",x"75",x"55",x"31",x"2d",x"51",x"55",x"75",x"71",x"71",x"75",x"51",x"30",x"51",x"55",x"75",x"51",x"6c",x"71",x"70",x"50",x"51",x"51",x"50",x"50",x"2d",x"04",x"04",x"08",x"08",x"51",x"b8",x"98",x"95",x"4d",x"2d",x"2d",x"0d",x"0d",x"0d",x"0d",x"2d",x"2d",x"2c",x"50",x"74",x"75",x"55",x"12",x"12",x"12",x"75",x"75",x"12",x"16",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"4d",x"71"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"05",x"09",x"29",x"88",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"ec",x"ec",x"cc",x"c8",x"a8",x"a8",x"c8",x"e8",x"e8",x"c8",x"a8",x"84",x"a8",x"c8",x"e8",x"49",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2e",x"32",x"32",x"4e",x"4e",x"2e",x"2e",x"2e",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"09",x"09",x"09",x"09",x"09",x"24",x"05",x"09",x"09",x"49",x"29",x"29",x"29",x"29",x"29",x"2d",x"32",x"4e",x"2e",x"32",x"32",x"32",x"2e",x"2d",x"54",x"55",x"51",x"55",x"51",x"31",x"31",x"31",x"30",x"30",x"11",x"11",x"11",x"12",x"12",x"11",x"11",x"12",x"12",x"12",x"75",x"b8",x"94",x"94",x"70",x"94",x"94",x"70",x"6c",x"4c",x"6c",x"4c",x"4c",x"70",x"70",x"70",x"70",x"70",x"6d",x"09",x"09",x"09",x"2d",x"75",x"94",x"70",x"70",x"71",x"4c",x"28",x"4c",x"70",x"75",x"94",x"94",x"94",x"95",x"95",x"95",x"72",x"6e",x"6d",x"6e",x"4d",x"4d",x"6d",x"49",x"05",x"29",x"4d",x"4d",x"49",x"4d",x"32",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"29",x"28",x"0d",x"09",x"09",x"28",x"28",x"0e",x"0d",x"09",x"09",x"2c",x"50",x"70",x"94",x"b4",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"99",x"b9",x"b9",x"b9",x"b9",x"95",x"71",x"4d",x"71",x"b5",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"2d",x"0d",x"09",x"09",x"09",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"55",x"75",x"51",x"2d",x"51",x"55",x"75",x"71",x"71",x"55",x"51",x"30",x"51",x"55",x"75",x"51",x"70",x"70",x"70",x"50",x"51",x"51",x"50",x"50",x"2c",x"08",x"04",x"08",x"08",x"2c",x"b8",x"b8",x"74",x"51",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"50",x"50",x"74",x"75",x"75",x"12",x"12",x"12",x"12",x"51",x"75",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"09",x"09",x"05",x"05",x"05",x"05",x"2d",x"95",x"b9"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"05",x"49",x"a8",x"e8",x"c8",x"a8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"ec",x"ec",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"cc",x"ec",x"ec",x"ec",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"ec",x"cc",x"c8",x"a8",x"c8",x"a8",x"cc",x"ec",x"ec",x"ec",x"cc",x"c8",x"a8",x"a8",x"e8",x"e8",x"c8",x"ec",x"c8",x"84",x"84",x"a8",x"e8",x"a8",x"29",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2e",x"32",x"32",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"25",x"05",x"09",x"09",x"09",x"09",x"24",x"25",x"09",x"29",x"4d",x"2d",x"49",x"49",x"29",x"2d",x"2d",x"2e",x"4e",x"2e",x"2e",x"2e",x"32",x"2e",x"2d",x"55",x"55",x"55",x"55",x"51",x"31",x"30",x"31",x"31",x"50",x"31",x"16",x"16",x"16",x"16",x"12",x"11",x"12",x"12",x"12",x"55",x"b8",x"b8",x"b8",x"94",x"70",x"4c",x"4c",x"70",x"71",x"4c",x"4c",x"4c",x"4c",x"70",x"70",x"70",x"70",x"71",x"09",x"0d",x"09",x"51",x"98",x"94",x"95",x"75",x"70",x"70",x"4c",x"28",x"4c",x"74",x"74",x"94",x"95",x"91",x"72",x"72",x"72",x"92",x"72",x"72",x"6d",x"4d",x"6d",x"4d",x"49",x"4d",x"4d",x"4d",x"49",x"52",x"3a",x"36",x"36",x"36",x"36",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"28",x"29",x"0d",x"09",x"09",x"28",x"28",x"0d",x"09",x"09",x"0d",x"0d",x"09",x"29",x"28",x"4c",x"4c",x"70",x"70",x"70",x"94",x"70",x"70",x"b5",x"b9",x"b9",x"b9",x"b9",x"95",x"75",x"4d",x"71",x"95",x"b9",x"b9",x"b9",x"b9",x"b9",x"b5",x"2d",x"0d",x"09",x"09",x"09",x"0d",x"31",x"55",x"56",x"36",x"12",x"12",x"16",x"55",x"75",x"55",x"2d",x"31",x"55",x"55",x"51",x"71",x"55",x"51",x"31",x"51",x"55",x"55",x"50",x"71",x"70",x"70",x"51",x"50",x"50",x"51",x"30",x"2c",x"08",x"04",x"08",x"08",x"2d",x"94",x"b8",x"74",x"94",x"2c",x"09",x"2d",x"2d",x"31",x"30",x"30",x"55",x"75",x"75",x"55",x"16",x"16",x"16",x"12",x"12",x"12",x"31",x"31",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"51",x"b9",x"b9",x"99"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"88",x"e8",x"c8",x"a8",x"88",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"c8",x"c8",x"c8",x"c8",x"cc",x"cc",x"ec",x"ec",x"e8",x"c8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a8",x"a8",x"a8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"ec",x"cc",x"c8",x"a8",x"a8",x"c8",x"e8",x"c8",x"e8",x"ec",x"a8",x"84",x"84",x"c8",x"e8",x"49",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2e",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"4e",x"2e",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"25",x"25",x"25",x"04",x"05",x"09",x"24",x"05",x"09",x"29",x"4d",x"2d",x"4d",x"49",x"2d",x"2d",x"2e",x"2e",x"2e",x"2e",x"2e",x"32",x"32",x"2d",x"4d",x"51",x"55",x"51",x"55",x"51",x"31",x"31",x"31",x"31",x"30",x"31",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"55",x"b8",x"b8",x"b9",x"b9",x"94",x"70",x"70",x"70",x"70",x"70",x"6c",x"4c",x"4c",x"70",x"70",x"70",x"70",x"70",x"09",x"09",x"09",x"71",x"b8",x"94",x"95",x"94",x"74",x"70",x"4c",x"28",x"4c",x"70",x"71",x"71",x"92",x"72",x"72",x"72",x"92",x"92",x"72",x"72",x"6e",x"6d",x"4d",x"4d",x"4d",x"6d",x"4d",x"4d",x"49",x"31",x"1a",x"36",x"3a",x"36",x"36",x"36",x"36",x"36",x"32",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0d",x"28",x"09",x"0d",x"09",x"09",x"28",x"28",x"0d",x"09",x"09",x"0d",x"0d",x"0d",x"09",x"29",x"2d",x"2d",x"2c",x"2d",x"29",x"2d",x"2d",x"4d",x"b8",x"b9",x"b5",x"b9",x"b9",x"b9",x"95",x"51",x"4d",x"95",x"b9",x"b9",x"b9",x"95",x"95",x"95",x"2d",x"09",x"0d",x"2d",x"31",x"51",x"55",x"55",x"75",x"75",x"55",x"35",x"12",x"11",x"75",x"55",x"31",x"30",x"55",x"55",x"55",x"71",x"55",x"31",x"31",x"51",x"55",x"55",x"50",x"71",x"70",x"70",x"51",x"51",x"50",x"4c",x"2d",x"2c",x"08",x"04",x"08",x"08",x"28",x"74",x"b8",x"74",x"98",x"2c",x"08",x"2c",x"2c",x"51",x"51",x"75",x"75",x"51",x"31",x"11",x"0e",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"09",x"09",x"05",x"05",x"09",x"09",x"05",x"4d",x"99",x"99",x"99"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"88",x"e8",x"c8",x"a8",x"84",x"a8",x"e8",x"e8",x"e8",x"c8",x"cc",x"ec",x"ec",x"ec",x"cc",x"ec",x"cc",x"cc",x"c8",x"cc",x"cc",x"ec",x"ec",x"ec",x"e8",x"c8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"a8",x"a4",x"a8",x"a8",x"a8",x"c8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"c8",x"a8",x"88",x"c8",x"c8",x"c8",x"c8",x"ec",x"c8",x"a4",x"84",x"a4",x"ec",x"68",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"32",x"32",x"32",x"32",x"2e",x"2e",x"32",x"2e",x"2e",x"2e",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"25",x"24",x"24",x"25",x"09",x"24",x"05",x"09",x"29",x"4e",x"4d",x"4d",x"4d",x"2d",x"4e",x"4e",x"2d",x"2d",x"2e",x"32",x"32",x"32",x"31",x"50",x"51",x"51",x"51",x"55",x"51",x"31",x"31",x"31",x"31",x"30",x"15",x"16",x"16",x"16",x"16",x"12",x"12",x"12",x"12",x"12",x"55",x"b9",x"b8",x"b9",x"b9",x"b8",x"95",x"95",x"90",x"70",x"70",x"70",x"70",x"4c",x"6c",x"91",x"94",x"74",x"94",x"0d",x"09",x"2d",x"75",x"98",x"94",x"99",x"94",x"94",x"75",x"70",x"4c",x"4c",x"50",x"71",x"72",x"72",x"72",x"92",x"92",x"92",x"92",x"72",x"72",x"72",x"6e",x"4d",x"4d",x"6d",x"6d",x"6e",x"4d",x"4d",x"31",x"16",x"16",x"36",x"36",x"36",x"36",x"3a",x"3a",x"36",x"36",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"28",x"0d",x"0d",x"09",x"09",x"08",x"28",x"09",x"09",x"09",x"0d",x"0d",x"2d",x"4d",x"4d",x"4d",x"2d",x"2d",x"09",x"09",x"09",x"05",x"29",x"b8",x"b4",x"b4",x"b5",x"b9",x"b9",x"95",x"71",x"4d",x"71",x"95",x"b5",x"95",x"95",x"75",x"71",x"09",x"09",x"2d",x"51",x"54",x"54",x"55",x"54",x"74",x"94",x"99",x"75",x"51",x"0d",x"75",x"55",x"30",x"30",x"51",x"55",x"55",x"55",x"55",x"31",x"2d",x"51",x"55",x"55",x"4c",x"71",x"74",x"70",x"51",x"51",x"4c",x"2c",x"2d",x"2c",x"28",x"04",x"08",x"08",x"08",x"50",x"dc",x"94",x"98",x"50",x"2c",x"2c",x"2c",x"51",x"75",x"75",x"51",x"2d",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"05",x"2d",x"75",x"79",x"79"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"cc",x"c8",x"a4",x"84",x"a4",x"c8",x"ec",x"e8",x"e8",x"c8",x"c8",x"cc",x"ec",x"ec",x"cc",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"ec",x"ec",x"e8",x"e8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"a8",x"a4",x"a8",x"a8",x"ec",x"c8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"c8",x"84",x"84",x"a8",x"a4",x"88",x"a8",x"c8",x"e8",x"ec",x"cc",x"cc",x"ec",x"ec",x"ec",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"c8",x"a8",x"88",x"a8",x"c8",x"c8",x"c8",x"e8",x"e8",x"c8",x"a8",x"a8",x"ec",x"88",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"52",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"24",x"25",x"24",x"05",x"09",x"29",x"52",x"4e",x"4d",x"4d",x"4d",x"4e",x"4e",x"2e",x"2e",x"32",x"52",x"2e",x"2d",x"51",x"50",x"51",x"51",x"51",x"51",x"51",x"30",x"31",x"31",x"30",x"30",x"15",x"16",x"16",x"16",x"16",x"12",x"11",x"12",x"12",x"12",x"32",x"95",x"d8",x"b9",x"b9",x"94",x"90",x"90",x"71",x"51",x"51",x"70",x"70",x"4c",x"6c",x"94",x"94",x"94",x"70",x"2d",x"09",x"51",x"94",x"98",x"95",x"94",x"94",x"94",x"70",x"70",x"4c",x"48",x"6d",x"92",x"92",x"72",x"72",x"92",x"92",x"72",x"72",x"92",x"6e",x"6e",x"6e",x"6e",x"6d",x"6d",x"4d",x"6d",x"6d",x"6d",x"31",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"0e",x"0d",x"2d",x"31",x"51",x"51",x"51",x"51",x"31",x"2d",x"28",x"0d",x"09",x"09",x"09",x"08",x"28",x"09",x"09",x"09",x"0d",x"2d",x"50",x"70",x"50",x"51",x"74",x"75",x"75",x"71",x"2d",x"09",x"29",x"b8",x"b4",x"94",x"b4",x"b9",x"b9",x"b9",x"75",x"4d",x"51",x"95",x"95",x"95",x"95",x"75",x"51",x"09",x"31",x"50",x"51",x"51",x"31",x"31",x"31",x"50",x"55",x"55",x"75",x"75",x"75",x"55",x"55",x"30",x"31",x"51",x"55",x"55",x"55",x"51",x"31",x"2d",x"51",x"55",x"55",x"4c",x"71",x"95",x"71",x"4c",x"2c",x"2c",x"2c",x"2c",x"2d",x"29",x"08",x"08",x"08",x"08",x"2c",x"dc",x"b8",x"75",x"51",x"4c",x"2c",x"2c",x"50",x"50",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"29",x"4d",x"09",x"05",x"05",x"4d",x"75",x"51",x"51"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"69",x"c8",x"c8",x"84",x"84",x"a8",x"ec",x"e8",x"e8",x"e8",x"c8",x"a8",x"c8",x"ec",x"ec",x"ec",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"e8",x"e8",x"c8",x"a8",x"88",x"84",x"84",x"88",x"88",x"84",x"a4",x"a4",x"a8",x"ec",x"c8",x"c8",x"cc",x"ec",x"ec",x"ec",x"ec",x"cc",x"ec",x"e8",x"e8",x"c8",x"a8",x"84",x"84",x"84",x"84",x"a8",x"c8",x"e8",x"ec",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a8",x"88",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"e8",x"c8",x"c8",x"e8",x"68",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"52",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"49",x"49",x"25",x"24",x"24",x"25",x"05",x"29",x"2d",x"4e",x"4e",x"4e",x"4e",x"52",x"52",x"52",x"32",x"32",x"32",x"2d",x"51",x"50",x"50",x"51",x"51",x"51",x"51",x"51",x"30",x"31",x"31",x"31",x"30",x"31",x"12",x"16",x"16",x"16",x"16",x"12",x"16",x"12",x"12",x"16",x"55",x"b9",x"b8",x"94",x"95",x"75",x"55",x"35",x"31",x"2d",x"4d",x"70",x"70",x"6c",x"94",x"98",x"94",x"94",x"51",x"09",x"71",x"98",x"94",x"95",x"94",x"95",x"98",x"74",x"70",x"71",x"4d",x"72",x"92",x"92",x"92",x"92",x"72",x"72",x"72",x"72",x"92",x"72",x"72",x"72",x"72",x"72",x"6e",x"6e",x"6d",x"6d",x"6d",x"32",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3a",x"32",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0d",x"09",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"12",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"2d",x"31",x"51",x"51",x"71",x"71",x"71",x"70",x"71",x"51",x"51",x"2c",x"0d",x"0d",x"09",x"09",x"09",x"28",x"09",x"09",x"09",x"0d",x"4c",x"50",x"50",x"50",x"50",x"70",x"74",x"95",x"95",x"75",x"4d",x"4d",x"b4",x"b9",x"b8",x"b8",x"b9",x"b9",x"95",x"75",x"51",x"4d",x"71",x"75",x"95",x"95",x"75",x"51",x"2d",x"31",x"50",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"51",x"55",x"75",x"75",x"75",x"55",x"31",x"2d",x"31",x"55",x"55",x"55",x"51",x"31",x"31",x"51",x"55",x"51",x"4c",x"70",x"94",x"50",x"2c",x"2c",x"2c",x"2c",x"2c",x"2c",x"2d",x"08",x"08",x"28",x"08",x"28",x"b8",x"b8",x"75",x"75",x"50",x"2c",x"2c",x"2d",x"09",x"09",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"09",x"4d",x"51",x"75",x"95",x"4d",x"2d",x"51",x"75",x"75",x"51",x"51"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"09",x"09",x"09",x"05",x"a8",x"c8",x"a4",x"84",x"a8",x"c8",x"ec",x"c8",x"c8",x"c8",x"c8",x"a8",x"c8",x"ec",x"ec",x"ec",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"ec",x"cc",x"ec",x"e8",x"c8",x"a4",x"88",x"a8",x"84",x"84",x"88",x"84",x"84",x"84",x"a8",x"ec",x"c8",x"c8",x"c8",x"ec",x"ec",x"ec",x"ec",x"cc",x"ec",x"c8",x"c8",x"c8",x"c8",x"84",x"84",x"84",x"84",x"a8",x"c8",x"c8",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"cc",x"ec",x"ec",x"ec",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"45",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"2e",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"2d",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"49",x"4d",x"4d",x"29",x"24",x"24",x"25",x"05",x"04",x"24",x"2d",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2d",x"11",x"51",x"50",x"51",x"51",x"51",x"51",x"50",x"51",x"51",x"30",x"31",x"31",x"31",x"30",x"2d",x"0d",x"0d",x"16",x"16",x"16",x"16",x"16",x"12",x"16",x"16",x"16",x"79",x"b4",x"70",x"75",x"36",x"16",x"16",x"0d",x"09",x"2d",x"95",x"70",x"4c",x"74",x"b8",x"94",x"95",x"70",x"09",x"71",x"98",x"95",x"95",x"94",x"94",x"94",x"74",x"71",x"71",x"72",x"92",x"92",x"72",x"72",x"92",x"72",x"72",x"72",x"92",x"92",x"72",x"72",x"92",x"92",x"92",x"92",x"6e",x"6d",x"6d",x"6d",x"32",x"1a",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"2d",x"31",x"0e",x"0e",x"0e",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"2d",x"71",x"95",x"94",x"94",x"75",x"70",x"71",x"70",x"71",x"70",x"70",x"4d",x"0d",x"0d",x"09",x"09",x"09",x"28",x"09",x"09",x"09",x"0d",x"2c",x"4c",x"2c",x"2c",x"4c",x"51",x"50",x"74",x"94",x"98",x"95",x"71",x"94",x"b9",x"b9",x"b9",x"b9",x"94",x"95",x"95",x"71",x"4d",x"51",x"71",x"95",x"95",x"75",x"51",x"54",x"31",x"51",x"51",x"55",x"75",x"75",x"75",x"51",x"30",x"30",x"51",x"55",x"75",x"79",x"75",x"51",x"2d",x"31",x"55",x"55",x"51",x"55",x"31",x"31",x"51",x"55",x"51",x"4c",x"70",x"94",x"71",x"51",x"2d",x"2d",x"2c",x"2c",x"2c",x"2d",x"08",x"08",x"28",x"08",x"28",x"94",x"dd",x"71",x"74",x"50",x"29",x"29",x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"51",x"95",x"bd",x"bd",x"bd",x"95",x"75",x"b9",x"b9",x"99",x"55",x"51"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"12",x"0d",x"0d",x"0d",x"0d",x"09",x"05",x"c8",x"c8",x"a4",x"a8",x"c8",x"ec",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"c8",x"ec",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"ec",x"c8",x"cc",x"e8",x"c8",x"a4",x"84",x"a4",x"a8",x"a8",x"84",x"84",x"84",x"a4",x"c8",x"ec",x"c8",x"a8",x"c8",x"cc",x"ec",x"c8",x"ec",x"ec",x"ec",x"c8",x"c8",x"c8",x"e8",x"c8",x"a8",x"a8",x"a8",x"cc",x"ec",x"c8",x"ec",x"ec",x"ec",x"c8",x"cc",x"ec",x"ec",x"c8",x"a8",x"c8",x"c8",x"c8",x"e8",x"e8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a4",x"a4",x"a4",x"c4",x"a4",x"c4",x"68",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"4e",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"2e",x"4e",x"4d",x"29",x"29",x"2d",x"29",x"49",x"4e",x"4d",x"4e",x"4e",x"29",x"24",x"24",x"25",x"09",x"05",x"24",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"51",x"50",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"2d",x"2d",x"30",x"30",x"0d",x"09",x"09",x"12",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"36",x"16",x"16",x"12",x"0d",x"0d",x"0d",x"09",x"09",x"95",x"94",x"4c",x"70",x"b9",x"95",x"94",x"90",x"2d",x"75",x"95",x"95",x"95",x"94",x"94",x"94",x"74",x"71",x"6d",x"6e",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"4d",x"6d",x"32",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"56",x"32",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"71",x"95",x"b9",x"b9",x"b9",x"b9",x"99",x"32",x"0d",x"0e",x"52",x"99",x"99",x"75",x"52",x"0e",x"0d",x"0d",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"2d",x"71",x"95",x"94",x"95",x"95",x"74",x"70",x"70",x"50",x"70",x"70",x"50",x"50",x"50",x"2d",x"0d",x"09",x"09",x"09",x"28",x"09",x"09",x"09",x"09",x"0c",x"2c",x"2c",x"2c",x"4c",x"50",x"70",x"74",x"94",x"98",x"98",x"95",x"94",x"b8",x"b8",x"94",x"94",x"70",x"70",x"70",x"51",x"4d",x"51",x"71",x"71",x"75",x"95",x"71",x"30",x"51",x"55",x"55",x"79",x"79",x"79",x"75",x"75",x"55",x"51",x"31",x"31",x"55",x"75",x"79",x"55",x"2c",x"31",x"55",x"55",x"51",x"55",x"31",x"31",x"51",x"55",x"51",x"4d",x"71",x"91",x"91",x"92",x"92",x"71",x"71",x"6d",x"4d",x"2c",x"08",x"09",x"09",x"09",x"05",x"51",x"d8",x"70",x"75",x"51",x"09",x"05",x"09",x"05",x"05",x"05",x"09",x"09",x"05",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"31",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"b9",x"99",x"75",x"75"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"09",x"05",x"a8",x"c8",x"c8",x"c8",x"e8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"a8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"ec",x"ec",x"ec",x"c8",x"c8",x"ec",x"c8",x"a4",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"a8",x"c8",x"e8",x"c8",x"a8",x"a8",x"cc",x"ec",x"e8",x"ec",x"e8",x"ec",x"c8",x"a8",x"a8",x"e8",x"e8",x"c8",x"c8",x"c8",x"cc",x"c8",x"c8",x"ec",x"ec",x"cc",x"c8",x"c8",x"ec",x"c8",x"c8",x"a8",x"a8",x"a8",x"c8",x"c8",x"ec",x"c8",x"a8",x"a8",x"88",x"88",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"68",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4d",x"4d",x"4d",x"29",x"4e",x"4e",x"4d",x"4d",x"4d",x"4d",x"24",x"25",x"05",x"09",x"05",x"20",x"0d",x"0e",x"09",x"29",x"09",x"09",x"05",x"05",x"05",x"09",x"31",x"50",x"51",x"51",x"50",x"51",x"51",x"51",x"31",x"30",x"2d",x"2d",x"30",x"30",x"0d",x"29",x"2d",x"56",x"3a",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"12",x"0d",x"09",x"09",x"09",x"09",x"0d",x"94",x"b8",x"4c",x"70",x"99",x"b8",x"94",x"70",x"51",x"71",x"95",x"94",x"95",x"94",x"95",x"98",x"74",x"71",x"4d",x"4d",x"6e",x"6e",x"72",x"72",x"92",x"92",x"92",x"92",x"72",x"72",x"92",x"92",x"92",x"92",x"72",x"6e",x"4d",x"4d",x"4d",x"6d",x"51",x"36",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"56",x"36",x"12",x"0e",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"51",x"75",x"99",x"b9",x"dd",x"bd",x"dd",x"dd",x"b9",x"51",x"0e",x"0e",x"52",x"b9",x"bd",x"b9",x"95",x"75",x"31",x"11",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"31",x"71",x"95",x"94",x"94",x"74",x"75",x"74",x"74",x"50",x"50",x"4c",x"50",x"50",x"50",x"2c",x"2c",x"0d",x"09",x"09",x"09",x"28",x"09",x"09",x"09",x"09",x"2c",x"2c",x"28",x"2c",x"4c",x"50",x"70",x"75",x"74",x"74",x"94",x"98",x"98",x"75",x"71",x"71",x"70",x"70",x"70",x"70",x"51",x"4c",x"4c",x"51",x"71",x"75",x"75",x"51",x"31",x"51",x"55",x"75",x"55",x"55",x"55",x"55",x"75",x"75",x"55",x"31",x"31",x"51",x"55",x"75",x"75",x"30",x"30",x"31",x"55",x"55",x"51",x"31",x"30",x"51",x"75",x"75",x"71",x"91",x"91",x"92",x"92",x"b2",x"92",x"91",x"6d",x"6d",x"4d",x"29",x"09",x"09",x"09",x"05",x"29",x"b8",x"94",x"74",x"55",x"2d",x"05",x"05",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"0d",x"09",x"55",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"12",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"12",x"12",x"11",x"11",x"11",x"11",x"12",x"31",x"29",x"05",x"88",x"c8",x"e8",x"c8",x"c8",x"c4",x"c8",x"c8",x"a4",x"a8",x"a8",x"c8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"c8",x"cc",x"c8",x"c8",x"ec",x"c8",x"a4",x"84",x"84",x"84",x"84",x"84",x"84",x"a8",x"c8",x"ec",x"e8",x"a8",x"a8",x"a8",x"c8",x"ec",x"e8",x"ec",x"e8",x"e8",x"c8",x"a8",x"a4",x"c4",x"c8",x"e8",x"e8",x"e8",x"c8",x"a8",x"a8",x"cc",x"ec",x"c8",x"a8",x"c8",x"e8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"ec",x"a8",x"a8",x"a8",x"a8",x"a8",x"a4",x"a4",x"a4",x"88",x"a8",x"a8",x"49",x"09",x"09",x"0d",x"09",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"2d",x"2e",x"32",x"32",x"32",x"32",x"32",x"52",x"4e",x"2e",x"2e",x"2e",x"2e",x"4e",x"2e",x"2d",x"4e",x"4e",x"4e",x"4d",x"4e",x"4d",x"4d",x"4d",x"4d",x"4d",x"24",x"25",x"25",x"29",x"29",x"24",x"32",x"36",x"2d",x"2e",x"2e",x"09",x"09",x"09",x"09",x"09",x"31",x"30",x"31",x"51",x"30",x"50",x"51",x"51",x"31",x"30",x"31",x"31",x"30",x"2c",x"2d",x"72",x"96",x"ba",x"ba",x"7a",x"36",x"16",x"16",x"16",x"16",x"16",x"16",x"11",x"0d",x"09",x"09",x"09",x"09",x"0d",x"0d",x"2d",x"b8",x"b8",x"6c",x"4c",x"94",x"b8",x"94",x"70",x"71",x"71",x"94",x"98",x"94",x"94",x"95",x"95",x"74",x"6d",x"49",x"49",x"49",x"4d",x"6d",x"6e",x"72",x"92",x"92",x"72",x"72",x"92",x"92",x"72",x"72",x"72",x"6e",x"4d",x"4d",x"4d",x"4d",x"6d",x"6d",x"32",x"16",x"16",x"16",x"16",x"16",x"36",x"36",x"36",x"36",x"36",x"36",x"56",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"31",x"99",x"dd",x"b9",x"b9",x"99",x"99",x"99",x"99",x"99",x"55",x"32",x"0e",x"52",x"99",x"b9",x"b9",x"b9",x"b9",x"95",x"32",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"31",x"95",x"b8",x"99",x"74",x"70",x"70",x"74",x"74",x"75",x"50",x"50",x"2c",x"2c",x"4d",x"4c",x"2c",x"2c",x"0d",x"09",x"09",x"09",x"28",x"08",x"09",x"09",x"28",x"4c",x"2c",x"2c",x"2c",x"4c",x"50",x"70",x"71",x"71",x"74",x"94",x"98",x"94",x"2d",x"29",x"4d",x"71",x"94",x"90",x"70",x"70",x"4c",x"48",x"4d",x"71",x"75",x"74",x"2d",x"31",x"51",x"55",x"55",x"31",x"2d",x"2d",x"31",x"55",x"75",x"55",x"51",x"31",x"30",x"51",x"55",x"75",x"50",x"30",x"31",x"55",x"55",x"51",x"30",x"30",x"51",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"6d",x"2d",x"0d",x"09",x"05",x"05",x"b8",x"b8",x"50",x"74",x"75",x"05",x"05",x"09",x"0d",x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"05",x"05",x"0d",x"0d",x"75",x"75",x"75",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"b9",x"b9",x"b9"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"12",x"11",x"11",x"12",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"31",x"ad",x"cc",x"a8",x"29",x"a8",x"c8",x"c4",x"c4",x"c4",x"c4",x"a4",x"a4",x"a8",x"a8",x"a8",x"c8",x"cc",x"ec",x"ec",x"cc",x"c8",x"ec",x"ec",x"ec",x"cc",x"cc",x"cc",x"c8",x"c8",x"e8",x"ec",x"c8",x"a8",x"a4",x"a4",x"a4",x"a8",x"c8",x"c8",x"ec",x"c8",x"c8",x"a4",x"a8",x"c8",x"c8",x"e8",x"e8",x"c8",x"e8",x"e8",x"cc",x"c8",x"a4",x"a4",x"a4",x"a8",x"c4",x"a4",x"a4",x"a8",x"c8",x"cc",x"c8",x"c8",x"a8",x"c8",x"e8",x"c8",x"a8",x"84",x"88",x"a8",x"a8",x"a8",x"c8",x"ec",x"c8",x"a8",x"a8",x"a8",x"a8",x"84",x"a8",x"a8",x"88",x"a8",x"c8",x"68",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"05",x"05",x"05",x"09",x"09",x"2d",x"4d",x"71",x"71",x"91",x"b5",x"b5",x"d5",x"d9",x"d9",x"d9",x"b5",x"4d",x"0e",x"32",x"32",x"32",x"32",x"32",x"32",x"2e",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"4e",x"4d",x"4d",x"4e",x"2d",x"4d",x"4d",x"4d",x"2d",x"00",x"91",x"48",x"91",x"b5",x"29",x"2e",x"32",x"29",x"2e",x"32",x"71",x"d9",x"d5",x"b5",x"b5",x"51",x"31",x"51",x"31",x"30",x"50",x"51",x"51",x"31",x"30",x"31",x"30",x"2c",x"75",x"da",x"df",x"ff",x"ff",x"ff",x"df",x"de",x"ba",x"56",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"94",x"b8",x"94",x"4c",x"4c",x"70",x"95",x"74",x"74",x"70",x"71",x"95",x"94",x"94",x"94",x"71",x"72",x"6e",x"6e",x"4d",x"49",x"49",x"49",x"4d",x"6d",x"6e",x"72",x"92",x"92",x"92",x"72",x"72",x"6e",x"6e",x"6e",x"4d",x"4d",x"4d",x"4d",x"6d",x"6d",x"52",x"3a",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"5a",x"36",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"31",x"75",x"b9",x"b9",x"99",x"99",x"99",x"99",x"95",x"95",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"52",x"12",x"12",x"12",x"0e",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"51",x"95",x"98",x"98",x"94",x"75",x"75",x"75",x"70",x"50",x"4c",x"4d",x"4c",x"2c",x"2c",x"4c",x"4c",x"2c",x"0d",x"0e",x"09",x"09",x"09",x"08",x"08",x"09",x"09",x"4c",x"4c",x"2c",x"2c",x"4c",x"4c",x"71",x"74",x"74",x"75",x"95",x"94",x"98",x"98",x"2d",x"09",x"09",x"2d",x"51",x"70",x"70",x"50",x"4c",x"4c",x"4c",x"71",x"75",x"51",x"31",x"31",x"51",x"31",x"0d",x"09",x"0d",x"09",x"0e",x"32",x"55",x"55",x"55",x"51",x"31",x"30",x"51",x"55",x"55",x"31",x"31",x"55",x"51",x"51",x"10",x"31",x"71",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"71",x"6d",x"4d",x"2d",x"09",x"05",x"71",x"b8",x"74",x"51",x"75",x"51",x"29",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"51",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"b9",x"b9",x"99",x"99"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"31",x"8d",x"ec",x"e8",x"ec",x"68",x"cc",x"c8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"a8",x"c8",x"cc",x"ec",x"ec",x"c8",x"c8",x"a8",x"c8",x"ec",x"ec",x"c8",x"c8",x"cc",x"c8",x"c8",x"e8",x"e8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"e8",x"c8",x"a4",x"a4",x"a8",x"c8",x"c8",x"c8",x"e8",x"c8",x"cc",x"c8",x"e8",x"c8",x"c8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"cc",x"e8",x"c8",x"c8",x"a8",x"c8",x"c8",x"e8",x"c8",x"a4",x"84",x"88",x"a8",x"a4",x"c8",x"c8",x"cc",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"a8",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"4d",x"4d",x"51",x"71",x"95",x"95",x"b5",x"d9",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"91",x"2e",x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"4e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"4e",x"2d",x"4d",x"4d",x"2d",x"4d",x"4d",x"4e",x"2d",x"00",x"d5",x"48",x"91",x"d9",x"29",x"2e",x"2d",x"2d",x"32",x"2e",x"96",x"fd",x"fd",x"fd",x"fd",x"51",x"31",x"51",x"31",x"31",x"51",x"51",x"51",x"30",x"30",x"2c",x"30",x"71",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ba",x"72",x"71",x"71",x"4d",x"4d",x"51",x"51",x"51",x"4d",x"4d",x"4d",x"4d",x"71",x"94",x"94",x"98",x"70",x"4c",x"4c",x"70",x"70",x"70",x"50",x"70",x"74",x"94",x"94",x"95",x"71",x"72",x"72",x"72",x"6e",x"6d",x"4d",x"49",x"49",x"4d",x"4d",x"6e",x"72",x"72",x"72",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"4d",x"6d",x"4d",x"4d",x"69",x"4e",x"36",x"36",x"36",x"36",x"36",x"3a",x"3a",x"36",x"36",x"36",x"36",x"5a",x"56",x"32",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"12",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0e",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"2d",x"75",x"99",x"95",x"95",x"79",x"75",x"75",x"75",x"75",x"99",x"dd",x"b9",x"b9",x"b9",x"b9",x"99",x"99",x"99",x"99",x"99",x"52",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"31",x"95",x"b8",x"98",x"95",x"94",x"95",x"95",x"95",x"74",x"50",x"4c",x"4d",x"4c",x"4c",x"2c",x"2c",x"2c",x"28",x"0d",x"0d",x"09",x"09",x"09",x"08",x"28",x"09",x"2d",x"50",x"50",x"4c",x"4c",x"50",x"50",x"70",x"74",x"74",x"95",x"95",x"98",x"98",x"98",x"2d",x"09",x"09",x"09",x"2d",x"71",x"70",x"50",x"70",x"4c",x"48",x"70",x"75",x"31",x"31",x"31",x"55",x"51",x"2d",x"09",x"09",x"09",x"0e",x"0e",x"31",x"55",x"55",x"55",x"31",x"2c",x"31",x"55",x"55",x"51",x"31",x"51",x"31",x"51",x"2c",x"51",x"92",x"92",x"92",x"92",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"91",x"91",x"8d",x"4d",x"09",x"05",x"29",x"b8",x"98",x"75",x"75",x"75",x"51",x"2d",x"2d",x"0d",x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"0d",x"2d",x"51",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"75"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"12",x"11",x"12",x"8d",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"a8",x"a8",x"a4",x"a4",x"a8",x"a8",x"a8",x"a8",x"c8",x"ec",x"ec",x"c8",x"a8",x"a8",x"a8",x"a8",x"c8",x"cc",x"c8",x"c8",x"cc",x"cc",x"c8",x"c8",x"c8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"c8",x"c4",x"a4",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a4",x"a4",x"a8",x"a8",x"c8",x"e8",x"e8",x"e8",x"c8",x"a8",x"a8",x"c8",x"e8",x"c8",x"a8",x"84",x"84",x"84",x"a4",x"a8",x"c8",x"ec",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"a8",x"a8",x"a8",x"49",x"09",x"09",x"09",x"09",x"4d",x"71",x"b1",x"d5",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"f9",x"6d",x"2e",x"32",x"32",x"32",x"32",x"2e",x"2e",x"4e",x"2e",x"4e",x"4e",x"4e",x"2e",x"4e",x"4e",x"4e",x"4d",x"4d",x"4d",x"4e",x"4e",x"4d",x"2d",x"24",x"d5",x"48",x"6d",x"da",x"0e",x"32",x"29",x"31",x"2e",x"0a",x"51",x"f9",x"fd",x"fd",x"fd",x"51",x"30",x"30",x"30",x"31",x"31",x"51",x"51",x"30",x"10",x"0c",x"51",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"d9",x"ba",x"b9",x"94",x"94",x"94",x"98",x"74",x"2c",x"28",x"4c",x"70",x"50",x"50",x"70",x"74",x"95",x"72",x"72",x"72",x"72",x"92",x"92",x"92",x"6e",x"6e",x"4d",x"49",x"49",x"4d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"4d",x"6d",x"4d",x"4d",x"69",x"6d",x"52",x"16",x"12",x"12",x"36",x"3a",x"3a",x"36",x"36",x"3a",x"36",x"5a",x"5a",x"36",x"12",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"31",x"2d",x"0d",x"0d",x"2d",x"75",x"75",x"51",x"55",x"55",x"51",x"51",x"51",x"55",x"99",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"99",x"95",x"75",x"31",x"0d",x"0e",x"0e",x"12",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"2d",x"95",x"b8",x"98",x"98",x"94",x"94",x"95",x"95",x"95",x"74",x"70",x"71",x"50",x"51",x"4c",x"2c",x"2c",x"2c",x"28",x"28",x"28",x"28",x"09",x"09",x"08",x"28",x"09",x"2d",x"50",x"50",x"50",x"50",x"70",x"70",x"50",x"70",x"75",x"95",x"94",x"98",x"98",x"94",x"09",x"09",x"09",x"0d",x"09",x"2d",x"90",x"50",x"71",x"4c",x"4c",x"74",x"74",x"0c",x"31",x"51",x"95",x"b9",x"75",x"2d",x"09",x"09",x"0d",x"0e",x"0e",x"31",x"55",x"55",x"31",x"2c",x"30",x"31",x"55",x"55",x"51",x"31",x"31",x"31",x"51",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"92",x"91",x"91",x"91",x"8d",x"4d",x"09",x"05",x"71",x"b9",x"94",x"51",x"51",x"78",x"95",x"75",x"51",x"2d",x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"29",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"55",x"51",x"51"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"12",x"11",x"51",x"c8",x"e8",x"e8",x"c8",x"cc",x"ec",x"e8",x"ec",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"ec",x"cc",x"a8",x"a8",x"a8",x"84",x"a8",x"c8",x"c8",x"c8",x"c8",x"cc",x"ec",x"c8",x"c8",x"c4",x"c8",x"c8",x"c8",x"e8",x"e8",x"c8",x"c8",x"c4",x"c4",x"a4",x"a4",x"a8",x"a8",x"c8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"c8",x"e8",x"c8",x"a8",x"a8",x"c8",x"c8",x"e8",x"c8",x"a8",x"84",x"84",x"84",x"a8",x"c8",x"ec",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"6d",x"91",x"b5",x"b5",x"d9",x"d9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"f9",x"d5",x"6d",x"0d",x"2e",x"32",x"32",x"32",x"2e",x"2e",x"4e",x"4e",x"4e",x"2e",x"4e",x"4e",x"4e",x"4e",x"4d",x"4e",x"4e",x"4e",x"2e",x"2d",x"91",x"24",x"f9",x"48",x"49",x"76",x"32",x"2e",x"29",x"32",x"2e",x"09",x"51",x"d9",x"fd",x"fd",x"fd",x"51",x"30",x"50",x"30",x"31",x"30",x"30",x"75",x"71",x"51",x"71",x"d6",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"b5",x"94",x"74",x"74",x"70",x"50",x"4c",x"4c",x"4c",x"4c",x"50",x"70",x"70",x"71",x"72",x"72",x"92",x"92",x"72",x"72",x"92",x"92",x"72",x"6e",x"6d",x"4d",x"49",x"4d",x"6d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"6d",x"4d",x"4d",x"6d",x"6d",x"4d",x"12",x"0e",x"0e",x"0e",x"12",x"36",x"36",x"36",x"36",x"36",x"32",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0d",x"0d",x"0d",x"12",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"0d",x"31",x"75",x"95",x"99",x"99",x"2d",x"51",x"99",x"99",x"75",x"51",x"51",x"51",x"51",x"51",x"75",x"75",x"99",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"99",x"31",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"75",x"b8",x"b8",x"98",x"98",x"94",x"94",x"95",x"95",x"95",x"71",x"50",x"4c",x"4c",x"4c",x"4c",x"2c",x"2c",x"2c",x"2c",x"2c",x"28",x"28",x"28",x"09",x"09",x"28",x"09",x"4d",x"70",x"50",x"51",x"50",x"50",x"71",x"71",x"70",x"75",x"75",x"94",x"b8",x"95",x"4d",x"09",x"09",x"09",x"0d",x"09",x"2d",x"94",x"70",x"70",x"4c",x"50",x"75",x"50",x"08",x"2c",x"94",x"99",x"b9",x"99",x"71",x"0d",x"09",x"0d",x"0e",x"0e",x"0e",x"31",x"51",x"51",x"31",x"2c",x"31",x"31",x"51",x"51",x"31",x"31",x"51",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"8d",x"6d",x"49",x"05",x"09",x"75",x"b8",x"98",x"74",x"54",x"51",x"51",x"51",x"51",x"70",x"75",x"95",x"75",x"95",x"4d",x"4d",x"51",x"75",x"75",x"79",x"99",x"b9",x"b9",x"b9",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"51",x"51",x"51"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"12",x"11",x"12",x"12",x"8d",x"e8",x"e8",x"c8",x"c8",x"c8",x"cc",x"c8",x"e8",x"c8",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"ec",x"c8",x"c8",x"a4",x"a8",x"84",x"84",x"a8",x"c8",x"c8",x"a8",x"c8",x"c8",x"e8",x"cc",x"c8",x"a4",x"c4",x"c4",x"c8",x"c8",x"c8",x"c4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"c8",x"e8",x"c8",x"c8",x"e8",x"c8",x"c8",x"e8",x"c8",x"a8",x"a4",x"a4",x"c8",x"e8",x"e8",x"c8",x"a8",x"a4",x"a8",x"a8",x"c8",x"e8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a4",x"a8",x"b1",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"f9",x"f9",x"f9",x"fe",x"fd",x"fd",x"b5",x"4d",x"2d",x"2e",x"2e",x"32",x"32",x"2e",x"4e",x"2e",x"2e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"2e",x"2d",x"71",x"91",x"44",x"f9",x"69",x"25",x"52",x"2e",x"4d",x"29",x"32",x"2e",x"29",x"4d",x"d9",x"fd",x"fd",x"fd",x"51",x"30",x"51",x"31",x"30",x"30",x"75",x"ba",x"ba",x"b5",x"d6",x"fa",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"d9",x"b9",x"95",x"95",x"95",x"95",x"71",x"4c",x"4c",x"4c",x"4c",x"50",x"71",x"72",x"72",x"72",x"92",x"92",x"72",x"72",x"72",x"92",x"92",x"72",x"6e",x"6d",x"49",x"49",x"4d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"4d",x"4d",x"6d",x"6d",x"4d",x"0d",x"0d",x"0d",x"0e",x"0e",x"12",x"32",x"32",x"12",x"12",x"12",x"11",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"0e",x"12",x"0d",x"09",x"0d",x"12",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"51",x"75",x"b9",x"b9",x"dd",x"bd",x"75",x"99",x"dd",x"b9",x"75",x"55",x"71",x"51",x"55",x"75",x"75",x"99",x"99",x"b9",x"b9",x"b9",x"b9",x"b9",x"99",x"95",x"99",x"b9",x"b9",x"75",x"32",x"12",x"0e",x"0e",x"0e",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"98",x"b8",x"98",x"98",x"98",x"98",x"95",x"95",x"74",x"75",x"71",x"50",x"4c",x"2c",x"4c",x"50",x"2c",x"2c",x"2c",x"50",x"2c",x"2c",x"2c",x"28",x"09",x"09",x"28",x"09",x"4c",x"70",x"70",x"71",x"50",x"50",x"75",x"75",x"74",x"75",x"94",x"94",x"94",x"51",x"09",x"09",x"09",x"09",x"0d",x"09",x"2d",x"94",x"70",x"70",x"50",x"70",x"75",x"50",x"0c",x"50",x"b4",x"98",x"99",x"b9",x"95",x"2d",x"09",x"0d",x"0e",x"0e",x"0e",x"0d",x"31",x"51",x"31",x"2d",x"2d",x"31",x"31",x"31",x"31",x"51",x"71",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"8d",x"6c",x"29",x"05",x"2d",x"95",x"b8",x"98",x"74",x"74",x"74",x"94",x"98",x"b8",x"b9",x"dd",x"bd",x"bd",x"75",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"b9",x"b9",x"99",x"99",x"79",x"99",x"99",x"99",x"55",x"2d",x"31",x"31"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"a8",x"e8",x"c8",x"c8",x"e8",x"e8",x"c8",x"c8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"cc",x"c8",x"ec",x"c8",x"a8",x"a4",x"84",x"84",x"a8",x"c8",x"e8",x"c8",x"a8",x"c8",x"e8",x"e8",x"cc",x"c8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"c8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"a8",x"a8",x"a4",x"a8",x"c8",x"c8",x"e8",x"ec",x"e8",x"c8",x"c8",x"ec",x"e8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a4",x"a8",x"d1",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"ff",x"fe",x"fe",x"f9",x"6d",x"29",x"0e",x"2e",x"32",x"2e",x"2e",x"2e",x"2e",x"4e",x"4e",x"4e",x"4e",x"4e",x"2e",x"32",x"32",x"2d",x"6d",x"f9",x"8d",x"49",x"f9",x"6d",x"05",x"29",x"29",x"49",x"29",x"52",x"52",x"29",x"4d",x"d9",x"fd",x"fd",x"fd",x"51",x"0c",x"31",x"31",x"2c",x"51",x"ff",x"ff",x"ff",x"fe",x"fa",x"fa",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fa",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"d9",x"95",x"4c",x"4c",x"4c",x"2c",x"4d",x"72",x"72",x"92",x"92",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"6e",x"6e",x"6e",x"6d",x"49",x"49",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"4d",x"4d",x"4d",x"6d",x"4d",x"2d",x"0d",x"0d",x"0e",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"0d",x"09",x"0d",x"12",x"12",x"12",x"12",x"0e",x"12",x"0d",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"31",x"75",x"99",x"b9",x"99",x"99",x"b9",x"b9",x"b9",x"b9",x"b9",x"99",x"79",x"75",x"75",x"75",x"75",x"95",x"99",x"99",x"b9",x"b9",x"b9",x"b9",x"99",x"99",x"75",x"55",x"55",x"75",x"99",x"b9",x"b9",x"55",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"95",x"98",x"98",x"98",x"98",x"98",x"94",x"75",x"70",x"70",x"71",x"74",x"70",x"71",x"51",x"50",x"4c",x"2c",x"2c",x"2c",x"4c",x"4d",x"50",x"4d",x"28",x"08",x"28",x"28",x"09",x"28",x"70",x"94",x"94",x"70",x"71",x"75",x"74",x"94",x"b8",x"b8",x"94",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"51",x"b8",x"94",x"74",x"70",x"70",x"74",x"30",x"0c",x"70",x"95",x"94",x"94",x"b8",x"95",x"51",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"2d",x"31",x"31",x"31",x"2c",x"2d",x"31",x"31",x"31",x"71",x"96",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"92",x"91",x"91",x"92",x"91",x"91",x"91",x"6d",x"68",x"09",x"09",x"0d",x"71",x"b8",x"dc",x"dc",x"dc",x"dc",x"b8",x"b9",x"b9",x"b9",x"b9",x"b9",x"75",x"75",x"99",x"99",x"99",x"99",x"75",x"75",x"55",x"79",x"99",x"99",x"79",x"79",x"99",x"99",x"79",x"51",x"2d",x"31",x"31"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"12",x"11",x"11",x"0e",x"11",x"11",x"11",x"11",x"0d",x"09",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"c8",x"a4",x"a8",x"a8",x"c8",x"e8",x"c8",x"c8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a4",x"a4",x"a4",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"c8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a4",x"cd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"f5",x"f9",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"da",x"b5",x"91",x"4d",x"09",x"0a",x"0e",x"2e",x"2e",x"2e",x"2e",x"2e",x"2e",x"0e",x"09",x"0d",x"29",x"71",x"d9",x"fd",x"49",x"69",x"fd",x"6d",x"05",x"25",x"25",x"29",x"24",x"29",x"2d",x"29",x"4d",x"d9",x"fd",x"fd",x"fd",x"51",x"30",x"31",x"30",x"30",x"ba",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fa",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"dd",x"b5",x"4c",x"4c",x"4c",x"6d",x"92",x"72",x"72",x"92",x"72",x"72",x"92",x"72",x"72",x"72",x"6e",x"6e",x"6e",x"6e",x"6d",x"4d",x"49",x"6d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"4d",x"4d",x"4d",x"6d",x"4d",x"4d",x"52",x"32",x"0d",x"0e",x"0d",x"0d",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"12",x"0d",x"09",x"0d",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"0d",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"0e",x"12",x"12",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"55",x"79",x"99",x"99",x"99",x"99",x"99",x"99",x"b9",x"99",x"b9",x"b9",x"99",x"99",x"b9",x"b9",x"b9",x"99",x"99",x"99",x"b9",x"b9",x"b9",x"b9",x"99",x"99",x"75",x"31",x"51",x"51",x"75",x"b9",x"b9",x"99",x"75",x"31",x"0e",x"0e",x"0e",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"94",x"98",x"98",x"98",x"98",x"98",x"94",x"94",x"74",x"74",x"74",x"74",x"75",x"75",x"70",x"4c",x"4c",x"4c",x"4c",x"2c",x"50",x"51",x"50",x"71",x"2c",x"08",x"28",x"28",x"09",x"08",x"28",x"4d",x"51",x"70",x"94",x"94",x"94",x"70",x"71",x"4d",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"75",x"b9",x"b9",x"b9",x"95",x"75",x"50",x"2c",x"2c",x"70",x"70",x"70",x"94",x"94",x"94",x"4d",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"31",x"31",x"31",x"2d",x"2d",x"31",x"31",x"51",x"92",x"96",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"6d",x"68",x"09",x"09",x"09",x"2d",x"2d",x"51",x"71",x"71",x"51",x"51",x"95",x"b9",x"99",x"99",x"79",x"75",x"79",x"79",x"99",x"99",x"75",x"55",x"51",x"31",x"55",x"99",x"99",x"75",x"79",x"99",x"79",x"99",x"75",x"2d",x"2d",x"2d"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"12",x"11",x"12",x"12",x"12",x"11",x"0d",x"0d",x"29",x"25",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"cc",x"ec",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"c8",x"c8",x"c8",x"ec",x"e8",x"c8",x"c4",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"cc",x"ec",x"ec",x"ec",x"cc",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a4",x"a4",x"a4",x"a4",x"c4",x"c8",x"c8",x"c8",x"c8",x"a4",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"84",x"ac",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"f5",x"f5",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"d5",x"91",x"4d",x"4d",x"4d",x"4d",x"4e",x"2e",x"2e",x"4d",x"4e",x"4d",x"4d",x"4d",x"25",x"91",x"fd",x"fd",x"28",x"6d",x"fd",x"6d",x"00",x"25",x"25",x"25",x"24",x"24",x"29",x"09",x"6d",x"f9",x"fd",x"fd",x"fd",x"51",x"2c",x"31",x"2c",x"71",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fa",x"d5",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"70",x"4c",x"71",x"72",x"92",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"4d",x"49",x"6d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"4d",x"4d",x"4d",x"4d",x"6d",x"b6",x"96",x"72",x"52",x"32",x"32",x"32",x"32",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"12",x"12",x"12",x"0e",x"0d",x"09",x"0d",x"12",x"0e",x"0d",x"11",x"12",x"0e",x"0d",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"0e",x"12",x"12",x"0e",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"75",x"75",x"75",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"99",x"99",x"b9",x"99",x"99",x"99",x"75",x"51",x"51",x"51",x"51",x"75",x"99",x"b9",x"b9",x"75",x"31",x"0e",x"52",x"51",x"2d",x"0d",x"0d",x"0d",x"2d",x"94",x"98",x"98",x"98",x"98",x"98",x"94",x"94",x"94",x"95",x"94",x"74",x"95",x"75",x"70",x"4c",x"50",x"50",x"50",x"4c",x"51",x"51",x"50",x"71",x"2c",x"08",x"28",x"28",x"09",x"08",x"04",x"09",x"2d",x"71",x"71",x"70",x"71",x"4d",x"29",x"09",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"72",x"ba",x"da",x"da",x"db",x"b6",x"95",x"54",x"2c",x"4d",x"95",x"71",x"70",x"70",x"70",x"70",x"4d",x"05",x"09",x"0d",x"0e",x"0e",x"0e",x"0e",x"0d",x"51",x"31",x"31",x"2c",x"31",x"31",x"51",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"92",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"71",x"91",x"6d",x"2d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"75",x"99",x"99",x"79",x"79",x"79",x"79",x"79",x"99",x"99",x"51",x"31",x"31",x"31",x"55",x"99",x"75",x"55",x"99",x"79",x"79",x"99",x"75",x"51",x"51",x"51"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"12",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"11",x"0d",x"09",x"25",x"88",x"c8",x"e8",x"c8",x"c8",x"c8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"ec",x"e8",x"e8",x"c8",x"c8",x"a4",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"ec",x"cc",x"c8",x"c8",x"c8",x"ec",x"ec",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"84",x"84",x"ac",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fa",x"fa",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"ff",x"fe",x"fd",x"f9",x"f9",x"f9",x"b5",x"91",x"8d",x"6d",x"6d",x"8d",x"91",x"b5",x"f9",x"f9",x"48",x"48",x"fd",x"fd",x"24",x"8d",x"fd",x"6d",x"04",x"25",x"25",x"25",x"24",x"29",x"25",x"05",x"71",x"fd",x"fd",x"fd",x"fd",x"51",x"2c",x"2c",x"51",x"ba",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fa",x"fe",x"fa",x"d5",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"95",x"71",x"72",x"92",x"72",x"72",x"72",x"72",x"72",x"72",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"49",x"6d",x"6d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"4d",x"4d",x"4d",x"49",x"6d",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"da",x"b6",x"96",x"72",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0e",x"12",x"0e",x"0d",x"12",x"12",x"0d",x"0e",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"0e",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0d",x"2d",x"55",x"95",x"99",x"99",x"99",x"b9",x"99",x"99",x"99",x"b9",x"b9",x"b9",x"99",x"99",x"99",x"99",x"b9",x"b9",x"b9",x"99",x"99",x"b9",x"75",x"75",x"79",x"99",x"75",x"31",x"31",x"51",x"51",x"99",x"b9",x"b9",x"b9",x"99",x"0e",x"79",x"bd",x"75",x"0d",x"09",x"09",x"2d",x"94",x"98",x"98",x"98",x"98",x"98",x"94",x"94",x"94",x"95",x"95",x"94",x"95",x"75",x"50",x"50",x"71",x"71",x"50",x"51",x"71",x"50",x"51",x"50",x"4c",x"2c",x"08",x"28",x"09",x"08",x"04",x"2d",x"51",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"92",x"db",x"ff",x"ff",x"ff",x"db",x"ff",x"b6",x"99",x"74",x"31",x"92",x"fb",x"b6",x"95",x"70",x"70",x"70",x"2d",x"05",x"05",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"31",x"31",x"31",x"2d",x"0c",x"31",x"4d",x"6d",x"6d",x"71",x"91",x"91",x"92",x"92",x"92",x"92",x"92",x"91",x"92",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"6d",x"4d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"51",x"79",x"75",x"79",x"75",x"75",x"79",x"79",x"75",x"75",x"75",x"51",x"2d",x"2d",x"51",x"95",x"99",x"75",x"55",x"99",x"75",x"75",x"75",x"99",x"99",x"95",x"95"),
(x"12",x"0d",x"0d",x"0d",x"0d",x"11",x"11",x"11",x"11",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"09",x"29",x"69",x"a8",x"c8",x"e8",x"e8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"c8",x"c8",x"cc",x"ec",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"a4",x"a4",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"c8",x"c8",x"a8",x"a8",x"a8",x"c8",x"c8",x"ec",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"a4",x"a4",x"a4",x"84",x"84",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"a8",x"84",x"a8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"ff",x"ff",x"fe",x"fd",x"fd",x"f9",x"f9",x"d9",x"d5",x"d5",x"d5",x"d9",x"f9",x"f9",x"f9",x"fd",x"6d",x"44",x"d5",x"fd",x"04",x"b1",x"fd",x"6d",x"24",x"49",x"25",x"24",x"25",x"25",x"01",x"25",x"b5",x"fd",x"fd",x"fd",x"fd",x"51",x"0c",x"2c",x"71",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fe",x"fa",x"d5",x"d5",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fd",x"b5",x"72",x"72",x"92",x"72",x"92",x"92",x"72",x"72",x"72",x"6e",x"4d",x"4d",x"4d",x"6d",x"6e",x"6e",x"6e",x"6e",x"6e",x"4d",x"6d",x"6d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"4d",x"4d",x"49",x"4d",x"d9",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"da",x"ba",x"ba",x"9a",x"96",x"96",x"76",x"52",x"52",x"32",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0e",x"12",x"0e",x"0e",x"12",x"12",x"0d",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"31",x"55",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"95",x"75",x"75",x"75",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"51",x"75",x"99",x"95",x"75",x"51",x"51",x"51",x"75",x"99",x"99",x"b9",x"b9",x"96",x"b9",x"dd",x"b9",x"71",x"4e",x"2e",x"51",x"b5",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"99",x"94",x"95",x"74",x"74",x"74",x"50",x"50",x"75",x"75",x"71",x"51",x"51",x"70",x"50",x"51",x"50",x"4c",x"2c",x"08",x"28",x"09",x"09",x"2c",x"71",x"95",x"71",x"4d",x"75",x"29",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"72",x"b6",x"db",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"b6",x"b9",x"74",x"51",x"b6",x"fb",x"db",x"ba",x"96",x"95",x"50",x"29",x"05",x"05",x"09",x"09",x"0d",x"0d",x"0d",x"0e",x"2e",x"31",x"31",x"2d",x"2d",x"51",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"91",x"91",x"91",x"92",x"92",x"92",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"71",x"91",x"6d",x"2d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"31",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"75",x"51",x"55",x"79",x"79",x"75",x"75",x"75",x"75",x"75",x"75"),
(x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"11",x"0d",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"25",x"89",x"c8",x"e8",x"e8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"c8",x"c8",x"a8",x"a8",x"c8",x"e8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"a8",x"a4",x"84",x"84",x"a4",x"a4",x"a8",x"ec",x"ec",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"a8",x"a4",x"84",x"a4",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"cc",x"cc",x"cc",x"cc",x"cc",x"a4",x"a8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fa",x"f5",x"f5",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"ff",x"fe",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"b1",x"48",x"8d",x"fd",x"04",x"b1",x"fd",x"6d",x"49",x"6d",x"49",x"00",x"25",x"25",x"25",x"6d",x"d9",x"fd",x"fd",x"fd",x"fe",x"51",x"0c",x"30",x"96",x"ff",x"ff",x"fe",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d5",x"d5",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"b6",x"92",x"72",x"72",x"72",x"92",x"92",x"72",x"72",x"72",x"6e",x"6d",x"4d",x"49",x"4d",x"6d",x"6e",x"6e",x"6e",x"6e",x"4d",x"6d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"6e",x"6e",x"6d",x"4d",x"4d",x"4d",x"4d",x"91",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"da",x"96",x"76",x"52",x"32",x"32",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"12",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"0d",x"0e",x"12",x"12",x"0e",x"12",x"11",x"0d",x"0d",x"0d",x"0e",x"0d",x"2d",x"51",x"75",x"99",x"b9",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"b9",x"99",x"75",x"75",x"55",x"55",x"55",x"75",x"95",x"99",x"99",x"99",x"99",x"99",x"75",x"51",x"51",x"75",x"95",x"95",x"75",x"51",x"75",x"99",x"99",x"b9",x"ba",x"ba",x"da",x"da",x"da",x"fa",x"d6",x"92",x"92",x"92",x"d5",x"da",x"da",x"da",x"da",x"d9",x"d9",x"b5",x"b5",x"b5",x"95",x"95",x"75",x"50",x"75",x"75",x"70",x"50",x"50",x"70",x"50",x"50",x"51",x"51",x"50",x"28",x"08",x"08",x"09",x"09",x"50",x"b8",x"94",x"94",x"94",x"b8",x"51",x"09",x"09",x"09",x"09",x"09",x"09",x"4d",x"db",x"ff",x"ff",x"ff",x"fb",x"fb",x"db",x"db",x"fb",x"96",x"95",x"94",x"75",x"b6",x"fb",x"db",x"db",x"db",x"b5",x"71",x"09",x"05",x"05",x"09",x"09",x"09",x"09",x"0d",x"0d",x"0e",x"31",x"31",x"51",x"51",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"71",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"71",x"91",x"91",x"4d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"2d",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"95",x"75",x"75",x"51",x"51",x"75",x"79",x"79",x"79",x"55",x"51",x"55",x"55",x"55"),
(x"11",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"09",x"09",x"05",x"05",x"05",x"05",x"69",x"c8",x"e8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"e8",x"c8",x"a8",x"a8",x"88",x"84",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"ec",x"ec",x"ec",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"84",x"84",x"84",x"84",x"84",x"a8",x"ec",x"cc",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"a8",x"a8",x"a8",x"a4",x"c8",x"f1",x"f0",x"f0",x"f0",x"f0",x"f0",x"cc",x"cc",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"f5",x"f0",x"f5",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"ff",x"fe",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"f9",x"69",x"24",x"f9",x"24",x"b1",x"fd",x"6d",x"69",x"d9",x"d9",x"04",x"69",x"91",x"91",x"d9",x"fd",x"fd",x"f9",x"fd",x"fd",x"51",x"0c",x"71",x"da",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d5",x"d5",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"92",x"6e",x"6e",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"6d",x"4d",x"49",x"4d",x"6e",x"6e",x"6e",x"6d",x"4d",x"6e",x"6e",x"6d",x"6e",x"6e",x"6d",x"6d",x"6e",x"6e",x"6d",x"4d",x"4d",x"4d",x"4d",x"6d",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"ba",x"96",x"76",x"52",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"11",x"12",x"0d",x"0e",x"0e",x"32",x"95",x"b9",x"2d",x"09",x"2d",x"75",x"99",x"99",x"99",x"b9",x"b9",x"b9",x"b9",x"99",x"99",x"99",x"99",x"99",x"b9",x"95",x"55",x"51",x"51",x"51",x"51",x"51",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"51",x"51",x"51",x"71",x"75",x"75",x"75",x"95",x"ba",x"d6",x"f6",x"f2",x"f2",x"f2",x"f6",x"f2",x"f2",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f2",x"f2",x"f2",x"f2",x"f2",x"f6",x"f6",x"f6",x"fa",x"da",x"b5",x"95",x"74",x"50",x"70",x"70",x"70",x"51",x"51",x"51",x"70",x"70",x"2c",x"08",x"08",x"09",x"09",x"95",x"b5",x"70",x"70",x"b4",x"94",x"71",x"09",x"09",x"09",x"05",x"09",x"92",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"db",x"fb",x"fb",x"b6",x"95",x"98",x"b9",x"b7",x"db",x"db",x"db",x"db",x"db",x"92",x"29",x"05",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"31",x"71",x"92",x"92",x"92",x"92",x"71",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"71",x"71",x"71",x"71",x"91",x"91",x"91",x"91",x"71",x"71",x"91",x"91",x"4d",x"2d",x"0d",x"0d",x"0e",x"0d",x"09",x"31",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"75",x"75",x"75",x"79",x"55",x"51",x"31",x"31",x"31"),
(x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"64",x"a8",x"e8",x"e8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"c8",x"a8",x"a8",x"88",x"84",x"84",x"c8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a4",x"a4",x"a4",x"a8",x"a8",x"c8",x"ec",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"a8",x"c8",x"c8",x"cc",x"c8",x"a4",x"a4",x"a4",x"a4",x"c8",x"ec",x"f0",x"f0",x"ec",x"f0",x"f0",x"cc",x"cc",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"ff",x"fe",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"91",x"24",x"8d",x"24",x"b1",x"fd",x"91",x"69",x"d9",x"fd",x"24",x"8d",x"d9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"51",x"2c",x"95",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d5",x"d5",x"f5",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"6e",x"4e",x"6e",x"6e",x"72",x"6e",x"72",x"72",x"72",x"72",x"92",x"92",x"72",x"6e",x"6d",x"49",x"4d",x"6e",x"6e",x"6e",x"6d",x"4d",x"6e",x"6e",x"6d",x"6d",x"6e",x"6d",x"6d",x"6e",x"6d",x"6d",x"6d",x"4d",x"4d",x"4d",x"49",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"da",x"ba",x"9a",x"96",x"76",x"52",x"32",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"32",x"95",x"b9",x"bd",x"75",x"51",x"75",x"99",x"99",x"99",x"b9",x"99",x"99",x"99",x"b9",x"b9",x"99",x"99",x"99",x"99",x"99",x"75",x"51",x"51",x"51",x"51",x"51",x"31",x"75",x"99",x"99",x"75",x"99",x"99",x"99",x"75",x"51",x"2d",x"51",x"51",x"51",x"95",x"da",x"f6",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ee",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"d6",x"b5",x"95",x"70",x"70",x"70",x"51",x"51",x"70",x"94",x"4c",x"28",x"09",x"08",x"08",x"51",x"94",x"95",x"4c",x"70",x"94",x"74",x"75",x"09",x"05",x"09",x"29",x"92",x"db",x"ff",x"ff",x"fb",x"fb",x"fb",x"db",x"db",x"db",x"db",x"fb",x"da",x"95",x"94",x"b9",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"72",x"09",x"05",x"09",x"09",x"0d",x"0d",x"09",x"09",x"09",x"09",x"71",x"91",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"91",x"91",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"6d",x"4d",x"2d",x"0e",x"0e",x"0d",x"2d",x"55",x"75",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"31",x"31",x"51",x"31",x"51",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"51",x"31",x"31"),
(x"0d",x"0d",x"09",x"09",x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"49",x"c8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"c8",x"88",x"84",x"84",x"84",x"a8",x"c8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"ec",x"cc",x"c8",x"c8",x"c8",x"ec",x"ec",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"c8",x"c8",x"ec",x"ec",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"c8",x"cc",x"ec",x"ec",x"ec",x"cc",x"a8",x"a8",x"a8",x"c8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"cc",x"f5",x"f0",x"ec",x"ec",x"f0",x"f1",x"f5",x"f9",x"f9",x"f9",x"f9",x"fd",x"f9",x"f6",x"fa",x"fe",x"fe",x"fe",x"fe",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"d9",x"49",x"24",x"20",x"b1",x"fd",x"91",x"49",x"b5",x"fd",x"24",x"91",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"51",x"51",x"ba",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d6",x"d5",x"d5",x"d5",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"d5",x"4d",x"4e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"72",x"72",x"72",x"72",x"72",x"6e",x"6e",x"4d",x"4d",x"6d",x"6e",x"6e",x"6e",x"4d",x"6d",x"6e",x"6d",x"6d",x"6e",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"4d",x"49",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"96",x"76",x"32",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"75",x"d9",x"b9",x"b9",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"75",x"75",x"99",x"b9",x"95",x"99",x"99",x"99",x"99",x"75",x"51",x"51",x"51",x"31",x"51",x"51",x"95",x"99",x"75",x"75",x"99",x"99",x"99",x"99",x"55",x"51",x"2d",x"2d",x"2d",x"b6",x"f6",x"ee",x"ea",x"ea",x"ea",x"ea",x"ee",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ee",x"f2",x"f6",x"b5",x"75",x"50",x"71",x"50",x"70",x"74",x"95",x"2c",x"08",x"09",x"08",x"28",x"74",x"94",x"75",x"4c",x"70",x"95",x"74",x"71",x"09",x"09",x"4d",x"92",x"db",x"ff",x"fb",x"fb",x"db",x"fb",x"fb",x"db",x"db",x"db",x"db",x"fb",x"da",x"95",x"94",x"d9",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"4d",x"05",x"09",x"09",x"0d",x"0d",x"09",x"05",x"0d",x"09",x"8d",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"71",x"71",x"71",x"71",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"0e",x"0d",x"0d",x"51",x"75",x"75",x"75",x"79",x"99",x"99",x"99",x"75",x"75",x"75",x"75",x"55",x"51",x"51",x"51",x"51",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"51",x"51"),
(x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"48",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"c8",x"a4",x"84",x"84",x"84",x"a4",x"c8",x"e8",x"c8",x"c8",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"c8",x"c8",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"c8",x"e8",x"e8",x"ec",x"e8",x"e8",x"c8",x"c8",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c8",x"cc",x"f0",x"f0",x"c8",x"ec",x"f0",x"f0",x"ec",x"cc",x"ec",x"cc",x"ec",x"ec",x"ec",x"cc",x"a8",x"88",x"a8",x"a8",x"a8",x"88",x"a8",x"cc",x"f1",x"ec",x"f0",x"ec",x"ec",x"c8",x"cc",x"f9",x"f9",x"f9",x"f9",x"fd",x"fa",x"fa",x"fe",x"ff",x"ff",x"fe",x"ff",x"ff",x"ff",x"fe",x"fa",x"fa",x"ff",x"ff",x"fa",x"fe",x"fe",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"b5",x"00",x"20",x"b5",x"fd",x"91",x"48",x"b5",x"dd",x"00",x"b1",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"75",x"71",x"da",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"da",x"d5",x"d5",x"d5",x"d1",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"b5",x"49",x"49",x"4d",x"4d",x"49",x"4d",x"4d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"4d",x"4d",x"6d",x"6e",x"6d",x"6e",x"4d",x"6d",x"6d",x"6d",x"4d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"6d",x"4d",x"4d",x"49",x"da",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"ba",x"96",x"72",x"32",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"12",x"12",x"0e",x"55",x"b9",x"b9",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"95",x"75",x"51",x"51",x"51",x"75",x"99",x"75",x"99",x"99",x"99",x"99",x"75",x"51",x"2d",x"2d",x"31",x"51",x"75",x"99",x"99",x"75",x"75",x"99",x"99",x"99",x"99",x"79",x"75",x"51",x"51",x"91",x"f6",x"ee",x"ea",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ee",x"ee",x"ee",x"f6",x"95",x"50",x"71",x"74",x"b4",x"94",x"2d",x"08",x"08",x"09",x"29",x"50",x"95",x"95",x"50",x"70",x"94",x"74",x"50",x"50",x"29",x"92",x"db",x"fb",x"fb",x"fb",x"ff",x"fb",x"fb",x"fb",x"db",x"db",x"db",x"db",x"db",x"fb",x"da",x"95",x"94",x"b9",x"ba",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b2",x"09",x"09",x"09",x"0d",x"0d",x"09",x"05",x"09",x"6d",x"91",x"91",x"91",x"91",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"92",x"91",x"91",x"91",x"91",x"91",x"91",x"71",x"71",x"91",x"71",x"71",x"71",x"71",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"4d",x"0e",x"0d",x"55",x"75",x"75",x"99",x"b9",x"99",x"99",x"b9",x"95",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75"),
(x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"09",x"05",x"05",x"09",x"29",x"88",x"c8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"c8",x"a4",x"84",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c4",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c4",x"c4",x"c4",x"e8",x"c8",x"c8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"cc",x"f0",x"f0",x"f0",x"a8",x"ec",x"f0",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"cc",x"a8",x"a8",x"a8",x"88",x"88",x"a8",x"ac",x"cc",x"ec",x"ec",x"f0",x"ec",x"ec",x"c8",x"d0",x"f9",x"fd",x"fd",x"f9",x"fd",x"fa",x"f5",x"f5",x"fa",x"fe",x"fe",x"fe",x"ff",x"fe",x"fe",x"fa",x"ff",x"ff",x"ff",x"ff",x"fe",x"fa",x"fa",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"fe",x"fd",x"f9",x"fd",x"fe",x"fe",x"fe",x"fd",x"f9",x"6d",x"8d",x"da",x"fe",x"b5",x"6d",x"b1",x"d9",x"00",x"d5",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"d9",x"ba",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"da",x"d5",x"d5",x"d5",x"d5",x"b1",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"d5",x"49",x"49",x"4d",x"49",x"49",x"49",x"4d",x"4d",x"6e",x"6e",x"6e",x"6e",x"6d",x"6e",x"6e",x"6d",x"49",x"6d",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"4d",x"49",x"49",x"b5",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"ba",x"9a",x"76",x"76",x"56",x"52",x"32",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"11",x"0e",x"32",x"75",x"b9",x"99",x"99",x"79",x"79",x"79",x"79",x"99",x"99",x"75",x"51",x"31",x"31",x"51",x"99",x"99",x"75",x"99",x"99",x"79",x"99",x"99",x"75",x"51",x"51",x"75",x"75",x"99",x"99",x"75",x"51",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"75",x"d6",x"f2",x"ee",x"ea",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"ee",x"f6",x"b5",x"74",x"74",x"74",x"70",x"4d",x"09",x"08",x"08",x"09",x"29",x"70",x"50",x"70",x"4c",x"4c",x"50",x"50",x"95",x"b5",x"92",x"db",x"ff",x"ff",x"fb",x"ff",x"ff",x"ff",x"fb",x"fb",x"db",x"db",x"db",x"fb",x"db",x"fb",x"fb",x"95",x"74",x"b8",x"b9",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"4d",x"09",x"09",x"0d",x"09",x"09",x"05",x"4d",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"92",x"91",x"92",x"92",x"91",x"91",x"91",x"91",x"91",x"91",x"71",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"0d",x"51",x"75",x"75",x"99",x"99",x"95",x"75",x"75",x"99",x"99",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"99",x"99",x"99",x"95",x"75",x"75",x"75",x"75"),
(x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"05",x"09",x"05",x"09",x"68",x"c4",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a4",x"a8",x"c8",x"ec",x"c8",x"c8",x"c4",x"a4",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"c8",x"a8",x"a4",x"84",x"88",x"88",x"84",x"a4",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"cc",x"f0",x"f1",x"cc",x"cc",x"a8",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"cc",x"cc",x"ac",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"ec",x"f0",x"ec",x"ec",x"f0",x"ec",x"f1",x"f9",x"f9",x"f9",x"f9",x"fd",x"fa",x"f1",x"ec",x"f4",x"fa",x"fe",x"fe",x"ff",x"fe",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fa",x"fa",x"f9",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"fe",x"f9",x"fd",x"f9",x"fa",x"ff",x"fe",x"da",x"b1",x"b1",x"b5",x"00",x"f9",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"da",x"d5",x"d5",x"d5",x"d5",x"d5",x"b1",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"d9",x"49",x"49",x"4d",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"4d",x"6d",x"6d",x"49",x"49",x"b5",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"b6",x"76",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"12",x"0e",x"51",x"75",x"99",x"79",x"75",x"79",x"79",x"79",x"79",x"99",x"99",x"75",x"31",x"31",x"51",x"75",x"99",x"75",x"55",x"79",x"79",x"99",x"79",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"51",x"51",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"79",x"95",x"f6",x"ee",x"ea",x"ea",x"ee",x"ee",x"ee",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ca",x"ca",x"ca",x"ee",x"ee",x"ee",x"f6",x"d5",x"94",x"94",x"70",x"2c",x"09",x"09",x"28",x"08",x"09",x"08",x"50",x"08",x"28",x"28",x"2c",x"4c",x"71",x"da",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"df",x"db",x"fb",x"fb",x"fb",x"fb",x"fb",x"db",x"db",x"db",x"95",x"74",x"b8",x"b9",x"db",x"db",x"db",x"db",x"db",x"db",x"d7",x"b6",x"92",x"09",x"09",x"0d",x"09",x"09",x"09",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"92",x"92",x"91",x"91",x"91",x"91",x"91",x"71",x"71",x"71",x"91",x"71",x"71",x"71",x"91",x"91",x"6d",x"71",x"71",x"71",x"6d",x"6d",x"6d",x"6d",x"2d",x"55",x"75",x"99",x"99",x"75",x"51",x"31",x"55",x"99",x"99",x"75",x"75",x"75",x"75",x"55",x"75",x"75",x"75",x"75",x"99",x"b9",x"b9",x"b9",x"b9",x"99",x"75",x"75",x"75",x"75"),
(x"09",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"09",x"49",x"a8",x"c4",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"c8",x"c8",x"c8",x"e8",x"c8",x"c4",x"c4",x"a4",x"a4",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c4",x"cc",x"d1",x"b5",x"b5",x"b9",x"b9",x"b5",x"b1",x"a4",x"84",x"ac",x"b5",x"b9",x"b1",x"ac",x"a4",x"c4",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"cc",x"f0",x"f0",x"ec",x"cc",x"ac",x"88",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"f0",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f1",x"f5",x"f9",x"fd",x"fa",x"fa",x"fa",x"f5",x"f9",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"ff",x"fa",x"fe",x"ff",x"ff",x"fa",x"ff",x"ff",x"ff",x"fa",x"d5",x"fa",x"fa",x"ff",x"fe",x"fe",x"fe",x"fe",x"da",x"91",x"48",x"fd",x"fe",x"fe",x"ff",x"ff",x"fe",x"fe",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"b1",x"d5",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"49",x"49",x"4d",x"49",x"49",x"4d",x"49",x"49",x"6d",x"6d",x"6d",x"6e",x"6d",x"6d",x"6d",x"6d",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"91",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"de",x"da",x"b6",x"76",x"32",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"0e",x"12",x"0e",x"31",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"95",x"75",x"75",x"99",x"99",x"75",x"55",x"55",x"99",x"79",x"99",x"75",x"75",x"75",x"75",x"79",x"95",x"75",x"75",x"51",x"51",x"55",x"75",x"99",x"79",x"79",x"79",x"99",x"79",x"99",x"ba",x"f2",x"ea",x"ea",x"ee",x"ee",x"ea",x"ca",x"ca",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ee",x"ee",x"ee",x"f6",x"f6",x"f2",x"f2",x"d6",x"92",x"09",x"09",x"28",x"08",x"09",x"09",x"4c",x"2c",x"2c",x"08",x"4d",x"b6",x"fb",x"fb",x"ff",x"ff",x"fb",x"ff",x"ff",x"fb",x"da",x"b6",x"d6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"d7",x"b5",x"94",x"94",x"b8",x"da",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"92",x"4d",x"09",x"0d",x"09",x"09",x"6d",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"92",x"91",x"91",x"91",x"91",x"71",x"71",x"71",x"91",x"71",x"71",x"71",x"71",x"71",x"71",x"71",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"55",x"75",x"99",x"75",x"31",x"31",x"31",x"75",x"99",x"79",x"75",x"55",x"75",x"55",x"75",x"75",x"55",x"75",x"99",x"99",x"79",x"75",x"75",x"79",x"99",x"99",x"75",x"75",x"75"),
(x"09",x"05",x"05",x"05",x"05",x"09",x"05",x"05",x"05",x"09",x"29",x"88",x"c8",x"a4",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"a4",x"a4",x"a4",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"b1",x"b5",x"b9",x"b9",x"b9",x"9d",x"9d",x"99",x"b1",x"84",x"80",x"ac",x"99",x"9d",x"b9",x"b5",x"b0",x"cc",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"f1",x"f0",x"cc",x"a8",x"88",x"a8",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"f1",x"f5",x"f9",x"f9",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"da",x"fe",x"ff",x"fa",x"fa",x"ff",x"ff",x"fe",x"d6",x"d5",x"fa",x"fe",x"ff",x"fa",x"ff",x"ff",x"fe",x"fe",x"b6",x"b1",x"f9",x"fa",x"da",x"d6",x"da",x"fa",x"fe",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d6",x"d6",x"fa",x"fa",x"fa",x"d5",x"d1",x"d5",x"d5",x"d5",x"d5",x"d5",x"b1",x"d5",x"f5",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fd",x"f9",x"4d",x"49",x"49",x"49",x"49",x"4d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"4d",x"6d",x"6d",x"49",x"91",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"9a",x"76",x"56",x"52",x"32",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"0e",x"0e",x"12",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"95",x"75",x"51",x"51",x"55",x"79",x"79",x"79",x"75",x"75",x"51",x"75",x"75",x"55",x"51",x"51",x"51",x"51",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"79",x"99",x"f6",x"f2",x"ea",x"ea",x"ee",x"ee",x"ea",x"ca",x"ca",x"ca",x"ea",x"ee",x"ee",x"ee",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"c9",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ee",x"ee",x"ee",x"f2",x"f2",x"ee",x"ee",x"f2",x"d2",x"72",x"2d",x"28",x"08",x"09",x"09",x"28",x"08",x"4c",x"6d",x"b6",x"fb",x"ff",x"fb",x"ff",x"db",x"fb",x"ff",x"ff",x"db",x"d6",x"b2",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"95",x"74",x"74",x"b8",x"ba",x"db",x"db",x"d6",x"da",x"db",x"d6",x"b6",x"92",x"6e",x"0d",x"0d",x"09",x"29",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"71",x"71",x"71",x"71",x"71",x"91",x"71",x"71",x"71",x"71",x"6d",x"71",x"6d",x"6d",x"6d",x"6d",x"71",x"6d",x"6d",x"51",x"79",x"99",x"55",x"31",x"31",x"51",x"75",x"79",x"75",x"55",x"55",x"75",x"55",x"75",x"75",x"55",x"75",x"99",x"75",x"55",x"51",x"51",x"55",x"75",x"99",x"99",x"75",x"75"),
(x"05",x"05",x"05",x"05",x"09",x"09",x"09",x"05",x"09",x"05",x"64",x"a8",x"a8",x"a4",x"a4",x"a4",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"d1",x"9d",x"9d",x"99",x"99",x"99",x"99",x"99",x"99",x"91",x"a8",x"84",x"90",x"99",x"99",x"99",x"99",x"99",x"b9",x"ac",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"ec",x"ec",x"cc",x"ac",x"88",x"88",x"a8",x"cc",x"f0",x"f0",x"f0",x"f0",x"cc",x"cc",x"cc",x"ac",x"cc",x"cc",x"d0",x"f0",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"f0",x"f0",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"f5",x"f5",x"f5",x"f5",x"fa",x"ff",x"fe",x"fe",x"fa",x"fa",x"fe",x"ff",x"ff",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"f9",x"f9",x"d5",x"d6",x"da",x"fe",x"fe",x"d6",x"fa",x"fe",x"ff",x"fa",x"d5",x"d5",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"fa",x"fe",x"fe",x"b1",x"b1",x"ad",x"88",x"a8",x"d1",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d6",x"d5",x"d5",x"d5",x"da",x"fa",x"fa",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d1",x"ad",x"d5",x"f5",x"f5",x"f5",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fd",x"fd",x"49",x"49",x"49",x"49",x"4d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"4d",x"6d",x"6d",x"49",x"6d",x"de",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"96",x"52",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"0e",x"11",x"12",x"12",x"12",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"75",x"79",x"79",x"79",x"75",x"51",x"51",x"51",x"51",x"31",x"31",x"51",x"51",x"75",x"75",x"99",x"b9",x"b9",x"b9",x"b9",x"99",x"99",x"b5",x"f6",x"ee",x"ee",x"ea",x"ee",x"ea",x"ca",x"ca",x"ca",x"ca",x"ea",x"ee",x"ee",x"ee",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"f6",x"91",x"28",x"08",x"09",x"09",x"28",x"08",x"71",x"fb",x"ff",x"ff",x"fb",x"fb",x"ff",x"da",x"fb",x"fb",x"ff",x"db",x"b6",x"b6",x"d6",x"db",x"fb",x"db",x"db",x"db",x"db",x"db",x"b6",x"b2",x"95",x"75",x"74",x"b8",x"b9",x"db",x"db",x"b6",x"d6",x"db",x"b6",x"b6",x"92",x"92",x"0d",x"09",x"09",x"4d",x"b1",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"71",x"71",x"71",x"71",x"71",x"91",x"91",x"6d",x"71",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"4d",x"75",x"79",x"55",x"31",x"51",x"99",x"75",x"75",x"51",x"51",x"55",x"55",x"55",x"75",x"55",x"75",x"99",x"79",x"55",x"31",x"51",x"51",x"31",x"51",x"75",x"99",x"75",x"55"),
(x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"09",x"05",x"29",x"84",x"a4",x"a8",x"a4",x"a8",x"a4",x"a8",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c8",x"b5",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"75",x"75",x"b5",x"b5",x"b5",x"99",x"99",x"79",x"79",x"99",x"99",x"99",x"ad",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c4",x"c8",x"c8",x"c8",x"c8",x"c8",x"ac",x"a8",x"88",x"88",x"a8",x"cc",x"f0",x"f0",x"f0",x"f0",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"f0",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"cc",x"f0",x"f0",x"cc",x"ac",x"ac",x"cc",x"cc",x"f0",x"f0",x"ec",x"f0",x"f0",x"f1",x"f5",x"fe",x"ff",x"fa",x"f1",x"f5",x"fe",x"ff",x"fa",x"ff",x"ff",x"fe",x"fa",x"f9",x"fa",x"fd",x"f9",x"d1",x"d6",x"fe",x"fa",x"d6",x"fe",x"ff",x"fe",x"f6",x"d5",x"d5",x"fa",x"fe",x"ff",x"fe",x"ff",x"ff",x"fe",x"fa",x"fa",x"fe",x"8d",x"64",x"64",x"64",x"84",x"88",x"b1",x"fa",x"fe",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d5",x"d5",x"d5",x"d5",x"d6",x"fa",x"fa",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"b1",x"ad",x"d5",x"f5",x"f5",x"f5",x"f9",x"fd",x"fd",x"fd",x"fe",x"fd",x"fd",x"fe",x"fe",x"fe",x"49",x"49",x"4d",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"4d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"de",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"de",x"de",x"ba",x"76",x"52",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"12",x"0e",x"51",x"75",x"75",x"75",x"75",x"99",x"75",x"75",x"75",x"75",x"75",x"55",x"51",x"51",x"31",x"51",x"51",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"51",x"51",x"51",x"51",x"51",x"55",x"75",x"99",x"99",x"99",x"95",x"99",x"99",x"99",x"b9",x"f6",x"f6",x"ee",x"ea",x"ea",x"ee",x"ea",x"ea",x"ca",x"ca",x"ca",x"ca",x"ee",x"ee",x"ee",x"ea",x"c9",x"ca",x"ee",x"ee",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ce",x"ca",x"c6",x"ca",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"f2",x"b1",x"29",x"09",x"09",x"28",x"72",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"fb",x"db",x"d7",x"db",x"db",x"fb",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"75",x"70",x"b8",x"b8",x"db",x"d7",x"d6",x"db",x"d7",x"b6",x"92",x"92",x"92",x"2d",x"09",x"2d",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"71",x"71",x"71",x"71",x"71",x"71",x"91",x"91",x"6d",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"75",x"79",x"95",x"75",x"75",x"75",x"55",x"51",x"31",x"51",x"55",x"55",x"55",x"55",x"55",x"75",x"79",x"75",x"31",x"31",x"31",x"31",x"31",x"31",x"75",x"99",x"75",x"55"),
(x"05",x"05",x"05",x"09",x"05",x"05",x"05",x"09",x"05",x"45",x"a4",x"a4",x"a4",x"a4",x"a8",x"a4",x"a4",x"a4",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a8",x"c8",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c8",x"b1",x"79",x"75",x"75",x"75",x"75",x"75",x"55",x"51",x"75",x"9d",x"b9",x"b9",x"99",x"99",x"99",x"79",x"75",x"75",x"59",x"91",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c4",x"c4",x"c8",x"c4",x"a4",x"a8",x"ac",x"ac",x"a8",x"a8",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"cc",x"a8",x"88",x"88",x"88",x"88",x"a8",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ac",x"f0",x"ec",x"ac",x"a8",x"a8",x"ac",x"ac",x"d0",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"fe",x"ff",x"fa",x"f0",x"f5",x"fe",x"fe",x"fa",x"ff",x"ff",x"ff",x"fa",x"f5",x"f9",x"f9",x"fd",x"d5",x"d6",x"da",x"da",x"d6",x"fe",x"ff",x"fe",x"d5",x"d5",x"f6",x"fa",x"fa",x"fe",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"b1",x"40",x"60",x"64",x"64",x"84",x"88",x"d1",x"fe",x"fe",x"fa",x"da",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d5",x"d1",x"d1",x"d5",x"d6",x"fa",x"fa",x"d5",x"d5",x"d5",x"d1",x"d1",x"d1",x"b1",x"b1",x"d5",x"f5",x"f5",x"f5",x"f9",x"f9",x"fd",x"fd",x"fe",x"fd",x"fd",x"fe",x"fe",x"d9",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"da",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"ba",x"76",x"56",x"52",x"32",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"12",x"31",x"75",x"75",x"75",x"95",x"99",x"99",x"99",x"75",x"75",x"75",x"75",x"75",x"51",x"51",x"51",x"51",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"51",x"51",x"75",x"75",x"75",x"99",x"99",x"95",x"75",x"55",x"55",x"75",x"b5",x"f6",x"f2",x"f2",x"ee",x"ea",x"ea",x"ee",x"ea",x"ea",x"ca",x"ca",x"ca",x"ca",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ea",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ee",x"f2",x"6d",x"09",x"09",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"ff",x"fb",x"fb",x"db",x"db",x"db",x"fb",x"fb",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ba",x"95",x"74",x"94",x"b8",x"da",x"db",x"da",x"db",x"b7",x"b6",x"92",x"92",x"92",x"4d",x"09",x"2d",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"8d",x"91",x"91",x"91",x"8d",x"8d",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"71",x"91",x"91",x"6d",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"51",x"55",x"75",x"75",x"75",x"51",x"51",x"31",x"31",x"51",x"55",x"55",x"55",x"55",x"55",x"75",x"75",x"75",x"31",x"31",x"31",x"31",x"31",x"51",x"75",x"79",x"55",x"55"),
(x"09",x"05",x"09",x"09",x"05",x"05",x"05",x"09",x"05",x"64",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"a4",x"a4",x"a8",x"a4",x"a4",x"a8",x"c8",x"c4",x"c4",x"c4",x"c8",x"c8",x"c4",x"c4",x"c4",x"ac",x"55",x"51",x"55",x"51",x"51",x"51",x"31",x"31",x"75",x"99",x"99",x"b9",x"b9",x"b9",x"b9",x"99",x"99",x"75",x"55",x"8c",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c4",x"c8",x"c4",x"a4",x"cc",x"f0",x"f0",x"cc",x"ec",x"ec",x"f0",x"ec",x"ec",x"f0",x"f0",x"cc",x"a8",x"88",x"88",x"88",x"88",x"a8",x"cc",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"ac",x"cc",x"ec",x"ac",x"88",x"88",x"a8",x"a8",x"cc",x"d0",x"ec",x"ec",x"ec",x"ec",x"c8",x"fa",x"fe",x"fa",x"f5",x"f9",x"fe",x"fa",x"fa",x"fe",x"ff",x"ff",x"fe",x"f9",x"f5",x"f5",x"fd",x"f9",x"b1",x"d1",x"d5",x"d5",x"fe",x"fe",x"fa",x"d1",x"d5",x"fa",x"f6",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"da",x"fe",x"fe",x"64",x"64",x"64",x"84",x"84",x"84",x"a8",x"d6",x"fe",x"fe",x"d6",x"d6",x"da",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d5",x"b1",x"d1",x"d5",x"d5",x"fa",x"d6",x"d5",x"d5",x"b1",x"b1",x"d1",x"b1",x"ad",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"fd",x"fe",x"fd",x"fd",x"fd",x"fd",x"fe",x"71",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"49",x"4d",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"b5",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"96",x"52",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"0e",x"55",x"75",x"75",x"99",x"b9",x"b9",x"99",x"b9",x"99",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"79",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"99",x"51",x"51",x"51",x"31",x"91",x"d2",x"f6",x"f2",x"ee",x"ee",x"ea",x"ee",x"ee",x"ea",x"ea",x"ca",x"ca",x"ca",x"ea",x"ca",x"ca",x"ca",x"f2",x"f6",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ee",x"ee",x"f2",x"f2",x"f6",x"f2",x"ea",x"ee",x"ea",x"ee",x"ea",x"ea",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"f2",x"b2",x"29",x"29",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"ff",x"fb",x"fb",x"fb",x"db",x"ff",x"db",x"db",x"db",x"fb",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"95",x"74",x"74",x"b8",x"da",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"4d",x"09",x"2d",x"8d",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"8d",x"6d",x"6d",x"8d",x"91",x"91",x"8d",x"91",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"91",x"71",x"6d",x"71",x"6d",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"4d",x"31",x"31",x"31",x"31",x"31",x"31",x"31",x"51",x"51",x"55",x"51",x"55",x"55",x"55",x"51",x"75",x"75",x"51",x"2d",x"31",x"31",x"31",x"75",x"79",x"75",x"51",x"55"),
(x"09",x"05",x"09",x"09",x"05",x"09",x"09",x"09",x"05",x"64",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a4",x"c8",x"c8",x"c4",x"c4",x"c8",x"cc",x"d1",x"b5",x"b5",x"c8",x"c8",x"b1",x"95",x"55",x"51",x"51",x"51",x"31",x"31",x"51",x"55",x"75",x"99",x"99",x"b9",x"b9",x"b9",x"b9",x"b9",x"b9",x"99",x"99",x"ac",x"c4",x"c4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c8",x"c4",x"c4",x"c4",x"c4",x"c8",x"cc",x"c8",x"a8",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"f0",x"f0",x"cc",x"cc",x"f0",x"f0",x"cc",x"ac",x"ac",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"ac",x"ac",x"cc",x"cc",x"cc",x"ac",x"88",x"a8",x"ac",x"d0",x"cc",x"cc",x"ec",x"cc",x"cc",x"fa",x"ff",x"fa",x"f5",x"fa",x"fe",x"fa",x"f9",x"fe",x"ff",x"ff",x"fe",x"f9",x"f5",x"f5",x"f9",x"fd",x"d5",x"d1",x"b1",x"b1",x"d5",x"d6",x"d5",x"b1",x"d5",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fe",x"ff",x"64",x"64",x"64",x"84",x"88",x"88",x"88",x"cd",x"fa",x"fe",x"fa",x"d6",x"d6",x"d6",x"da",x"fa",x"fa",x"fa",x"fa",x"fa",x"da",x"d6",x"d6",x"d5",x"b1",x"b1",x"d5",x"d5",x"fa",x"d6",x"d5",x"d1",x"d1",x"b1",x"ad",x"b1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"b9",x"49",x"49",x"6d",x"6d",x"4d",x"49",x"49",x"4d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"4d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"6d",x"da",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"ba",x"96",x"76",x"32",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"12",x"12",x"32",x"75",x"75",x"99",x"99",x"75",x"55",x"55",x"99",x"99",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"b9",x"b9",x"b9",x"99",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"95",x"51",x"31",x"51",x"51",x"d2",x"f2",x"f2",x"ee",x"ee",x"ee",x"ea",x"ee",x"ee",x"ee",x"ea",x"c9",x"c9",x"ca",x"ca",x"ca",x"ca",x"f2",x"f2",x"f2",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"f2",x"f2",x"ee",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"8d",x"52",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"df",x"df",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"95",x"54",x"70",x"b8",x"b6",x"b6",x"b7",x"b6",x"b6",x"92",x"92",x"92",x"8e",x"6d",x"29",x"29",x"6d",x"6d",x"8d",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"6d",x"6d",x"6d",x"8d",x"8d",x"91",x"8d",x"91",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"31",x"2d",x"2d",x"31",x"31",x"51",x"51",x"55",x"51",x"51",x"51",x"51",x"55",x"51",x"51",x"75",x"75",x"75",x"75",x"75",x"75",x"79",x"75",x"51",x"51",x"55"),
(x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"64",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c8",x"e4",x"c8",x"c8",x"ad",x"b5",x"b9",x"9d",x"bd",x"b1",x"b1",x"b9",x"99",x"55",x"51",x"51",x"51",x"51",x"51",x"55",x"75",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"b0",x"c8",x"c8",x"c4",x"c4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c4",x"c4",x"c4",x"c4",x"c8",x"ec",x"cc",x"cc",x"c8",x"f0",x"f0",x"cc",x"cc",x"d0",x"f0",x"ec",x"ec",x"f0",x"cc",x"cc",x"cc",x"f0",x"f0",x"cc",x"cc",x"cc",x"d0",x"cc",x"cc",x"a8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"ac",x"ac",x"cc",x"cc",x"cc",x"cc",x"ac",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"f5",x"fa",x"fa",x"f5",x"f5",x"fa",x"fa",x"f5",x"fa",x"fe",x"ff",x"fa",x"f5",x"f5",x"f5",x"f9",x"fd",x"f9",x"d1",x"b1",x"b1",x"d5",x"d1",x"b1",x"ad",x"d5",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"88",x"64",x"64",x"84",x"88",x"88",x"88",x"a8",x"d1",x"fe",x"fe",x"f6",x"d5",x"d5",x"d5",x"d6",x"d6",x"da",x"d6",x"d6",x"d5",x"d5",x"d5",x"d5",x"b1",x"b1",x"d1",x"d5",x"d5",x"d5",x"d5",x"d1",x"d1",x"b1",x"ad",x"d1",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"fe",x"fd",x"fd",x"fd",x"fe",x"fd",x"71",x"49",x"6d",x"6d",x"6e",x"6d",x"49",x"49",x"49",x"4d",x"49",x"29",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"4d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"b6",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"96",x"56",x"52",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"12",x"51",x"75",x"95",x"99",x"75",x"51",x"31",x"31",x"79",x"99",x"75",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"99",x"b9",x"b9",x"b9",x"99",x"95",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"75",x"31",x"31",x"31",x"51",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ee",x"ea",x"ea",x"ee",x"ea",x"c9",x"ca",x"ca",x"ca",x"ee",x"f2",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"f2",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c9",x"ea",x"ea",x"ea",x"ea",x"ee",x"d2",x"b6",x"ff",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"db",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"d6",x"95",x"54",x"50",x"b8",x"b5",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6e",x"6d",x"6d",x"4d",x"48",x"48",x"6d",x"6d",x"91",x"91",x"91",x"91",x"91",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"91",x"8d",x"8d",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"4d",x"51",x"31",x"31",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"55",x"51",x"31",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"31",x"51",x"55"),
(x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"64",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c8",x"c4",x"c4",x"c4",x"c8",x"c8",x"c4",x"c4",x"c4",x"ad",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"75",x"55",x"55",x"55",x"75",x"75",x"95",x"99",x"b9",x"99",x"99",x"99",x"99",x"75",x"51",x"51",x"75",x"99",x"99",x"b5",x"cd",x"c4",x"c4",x"c4",x"c4",x"c4",x"c8",x"c8",x"c4",x"c4",x"c4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c4",x"c4",x"c4",x"c4",x"cc",x"f0",x"cc",x"cc",x"f0",x"cc",x"ac",x"a8",x"ac",x"cc",x"f0",x"ec",x"ec",x"f0",x"cc",x"ac",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"a8",x"a8",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"a8",x"a8",x"cc",x"cc",x"d0",x"f0",x"d0",x"d0",x"ac",x"cc",x"ec",x"cc",x"ec",x"f0",x"f0",x"f0",x"f5",x"f5",x"f5",x"f9",x"f5",x"f1",x"f5",x"fa",x"fa",x"fa",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"d5",x"b1",x"d6",x"fa",x"d6",x"b1",x"8d",x"d5",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"fa",x"fa",x"fa",x"fa",x"fa",x"d6",x"b1",x"64",x"64",x"84",x"84",x"88",x"a8",x"a8",x"ad",x"fa",x"fe",x"fa",x"b5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"b1",x"b1",x"b1",x"d5",x"d5",x"d5",x"d1",x"d1",x"b1",x"b1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"fe",x"fe",x"fd",x"fe",x"fe",x"d9",x"49",x"4d",x"6e",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"4d",x"49",x"29",x"29",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"49",x"4d",x"49",x"91",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ba",x"76",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"0e",x"75",x"75",x"99",x"75",x"51",x"31",x"31",x"31",x"99",x"99",x"75",x"75",x"75",x"75",x"55",x"75",x"75",x"75",x"99",x"99",x"95",x"75",x"75",x"75",x"79",x"99",x"99",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"99",x"51",x"2d",x"2d",x"51",x"d2",x"ee",x"ea",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"ee",x"ee",x"ea",x"c9",x"ca",x"ca",x"f2",x"f2",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"c9",x"c9",x"ca",x"ea",x"ea",x"ea",x"f2",x"fb",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"da",x"b6",x"92",x"fa",x"fa",x"fa",x"f6",x"f6",x"f6",x"fa",x"fb",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"95",x"54",x"51",x"b8",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"6e",x"91",x"b1",x"8d",x"48",x"48",x"48",x"6d",x"8d",x"91",x"91",x"91",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"8d",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"4d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"51",x"51",x"55",x"55",x"51",x"51",x"31",x"31",x"51",x"55"),
(x"b5",x"b5",x"b5",x"b5",x"b5",x"b5",x"b5",x"b5",x"b5",x"a8",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"8c",x"75",x"79",x"79",x"79",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"31",x"51",x"51",x"55",x"99",x"99",x"b5",x"b1",x"c8",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c8",x"c8",x"c8",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"a4",x"c8",x"f0",x"f0",x"cc",x"cc",x"f0",x"ac",x"a8",x"88",x"a8",x"cc",x"cc",x"cc",x"cc",x"ec",x"cc",x"ac",x"a8",x"a8",x"ac",x"ac",x"ac",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"ec",x"ec",x"cc",x"cc",x"ec",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"ac",x"ac",x"cc",x"ac",x"ac",x"cc",x"cc",x"cc",x"ec",x"f0",x"f1",x"ac",x"cc",x"cc",x"f1",x"f1",x"f9",x"fa",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"d5",x"d1",x"fa",x"fe",x"fa",x"d1",x"ad",x"d5",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fa",x"fa",x"fa",x"fa",x"d1",x"fa",x"88",x"60",x"84",x"84",x"88",x"88",x"ad",x"a8",x"d1",x"fa",x"fe",x"d6",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d1",x"b1",x"b1",x"b1",x"d1",x"d1",x"d1",x"b1",x"b1",x"b1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"fe",x"fe",x"fd",x"fd",x"fd",x"b5",x"49",x"6d",x"6e",x"6d",x"6d",x"6e",x"6d",x"49",x"29",x"49",x"49",x"29",x"25",x"29",x"49",x"6d",x"6d",x"6d",x"6d",x"4d",x"6d",x"6d",x"6d",x"4d",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"4d",x"49",x"4d",x"b6",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"de",x"ba",x"9a",x"76",x"56",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0e",x"12",x"12",x"12",x"55",x"75",x"99",x"75",x"2d",x"2d",x"51",x"75",x"79",x"75",x"55",x"51",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"75",x"75",x"51",x"51",x"51",x"55",x"95",x"99",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"95",x"75",x"75",x"75",x"f2",x"ee",x"ea",x"ea",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"c9",x"ca",x"ca",x"f2",x"f2",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"c9",x"ca",x"ca",x"c9",x"ca",x"ca",x"c9",x"ca",x"ea",x"ea",x"ea",x"ee",x"fa",x"fb",x"fa",x"f6",x"f6",x"f6",x"f6",x"f6",x"d6",x"d6",x"f6",x"f2",x"f2",x"ee",x"ee",x"ee",x"f2",x"f6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ba",x"75",x"54",x"74",x"b8",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"91",x"91",x"8d",x"48",x"48",x"48",x"48",x"6d",x"6d",x"91",x"91",x"91",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"8d",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"31",x"31",x"51",x"51",x"31",x"2d",x"31",x"31",x"51",x"51"),
(x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"cd",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"91",x"55",x"55",x"75",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"b9",x"b9",x"99",x"99",x"b9",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"99",x"75",x"2d",x"2d",x"2d",x"31",x"75",x"99",x"99",x"99",x"b1",x"c8",x"c4",x"c8",x"ac",x"c8",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"a4",x"a4",x"ec",x"f0",x"cc",x"cc",x"f0",x"d0",x"a8",x"88",x"a8",x"ac",x"cc",x"cc",x"a8",x"cc",x"ec",x"ec",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"cc",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"ec",x"ec",x"cc",x"ec",x"f0",x"f1",x"a8",x"88",x"a8",x"cc",x"f1",x"f5",x"f9",x"f5",x"f5",x"d5",x"d5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"d5",x"f5",x"fa",x"fa",x"d1",x"b1",x"d5",x"fa",x"fe",x"fe",x"ff",x"ff",x"fe",x"ff",x"fa",x"fa",x"fa",x"fa",x"d1",x"fe",x"b1",x"64",x"64",x"84",x"88",x"88",x"a9",x"a8",x"ad",x"fa",x"fe",x"d6",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"b1",x"b1",x"ad",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"d5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"fd",x"fe",x"fe",x"fd",x"f9",x"91",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"25",x"49",x"49",x"29",x"29",x"29",x"49",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"6d",x"4d",x"4d",x"6d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"91",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ba",x"76",x"52",x"32",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"12",x"55",x"75",x"99",x"75",x"31",x"51",x"75",x"75",x"75",x"51",x"51",x"51",x"75",x"75",x"75",x"75",x"75",x"99",x"79",x"55",x"51",x"51",x"31",x"31",x"31",x"75",x"99",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"75",x"95",x"99",x"75",x"79",x"b5",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"ca",x"ca",x"ca",x"ee",x"f2",x"ca",x"ca",x"ea",x"ea",x"ca",x"ee",x"ea",x"ca",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"c9",x"ca",x"ca",x"c9",x"ca",x"ca",x"ca",x"c5",x"c9",x"e9",x"ea",x"ee",x"f6",x"fa",x"f6",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f6",x"f2",x"f2",x"ee",x"e9",x"c5",x"c5",x"e9",x"f6",x"fa",x"db",x"db",x"db",x"b6",x"b6",x"db",x"db",x"ba",x"95",x"54",x"50",x"94",x"b8",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"8d",x"91",x"91",x"8d",x"6d",x"48",x"48",x"48",x"48",x"6d",x"6d",x"91",x"91",x"91",x"8d",x"6d",x"6d",x"6d",x"6d",x"91",x"8d",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"48",x"4d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"31",x"31",x"51",x"51",x"51"),
(x"f9",x"f9",x"fd",x"fd",x"f9",x"f9",x"f9",x"fd",x"fd",x"d1",x"a4",x"84",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"a8",x"71",x"55",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"b9",x"b9",x"99",x"79",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"75",x"79",x"75",x"51",x"2d",x"2d",x"2d",x"51",x"75",x"99",x"99",x"99",x"b5",x"c4",x"b1",x"9d",x"b5",x"c8",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"a4",x"a4",x"a4",x"a4",x"a4",x"f0",x"f0",x"cc",x"cc",x"f1",x"cc",x"88",x"88",x"ac",x"cc",x"cc",x"ac",x"a8",x"cc",x"ec",x"ec",x"cc",x"cc",x"ac",x"ac",x"a8",x"a8",x"a8",x"ac",x"ac",x"cc",x"cc",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"cc",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"cc",x"ec",x"ec",x"cc",x"cc",x"f0",x"ec",x"cc",x"88",x"88",x"ac",x"cc",x"d1",x"d5",x"f5",x"fa",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"d5",x"b1",x"d1",x"b1",x"b1",x"d5",x"fa",x"fa",x"fa",x"ff",x"fa",x"fe",x"ff",x"fa",x"fa",x"fa",x"fa",x"b1",x"d5",x"fa",x"ad",x"64",x"64",x"88",x"88",x"a8",x"a8",x"ad",x"f6",x"fe",x"d5",x"b1",x"d1",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d1",x"b1",x"ad",x"b1",x"b1",x"ad",x"ad",x"b1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"fd",x"fd",x"fe",x"fe",x"d9",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"6d",x"4d",x"4d",x"6d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"4d",x"49",x"49",x"4d",x"49",x"4d",x"49",x"6d",x"da",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"96",x"56",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"12",x"31",x"55",x"51",x"75",x"95",x"75",x"79",x"75",x"75",x"51",x"31",x"51",x"51",x"55",x"55",x"55",x"75",x"75",x"79",x"75",x"51",x"31",x"31",x"31",x"31",x"31",x"55",x"79",x"75",x"55",x"55",x"55",x"55",x"75",x"51",x"31",x"51",x"55",x"55",x"35",x"51",x"b1",x"ee",x"ee",x"c9",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"c9",x"ca",x"ce",x"f2",x"f2",x"ca",x"ca",x"ca",x"ee",x"f2",x"ee",x"c9",x"ca",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"ce",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c5",x"c5",x"ee",x"f2",x"f6",x"fa",x"f6",x"f6",x"f2",x"ca",x"c9",x"e9",x"ea",x"ea",x"ee",x"f2",x"f2",x"ee",x"ea",x"c5",x"c5",x"c5",x"ee",x"f6",x"db",x"db",x"b6",x"6e",x"6d",x"b2",x"b6",x"95",x"74",x"50",x"74",x"b8",x"b9",x"92",x"92",x"92",x"b6",x"92",x"92",x"92",x"91",x"91",x"91",x"91",x"91",x"91",x"6d",x"48",x"48",x"48",x"48",x"48",x"6d",x"91",x"91",x"8d",x"8d",x"6d",x"8d",x"8d",x"91",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"48",x"48",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"48",x"48",x"4d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"31",x"31",x"51",x"51",x"51",x"51",x"51"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"a8",x"84",x"84",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c8",x"ad",x"75",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"75",x"55",x"75",x"75",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"51",x"75",x"75",x"75",x"51",x"51",x"2d",x"31",x"75",x"99",x"99",x"99",x"99",x"b1",x"95",x"7d",x"99",x"b1",x"c4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c8",x"cc",x"cc",x"cc",x"f0",x"cc",x"ac",x"ac",x"cc",x"cc",x"cc",x"a8",x"a8",x"cc",x"ec",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"f0",x"f0",x"f0",x"d0",x"d0",x"f0",x"f0",x"f0",x"f0",x"cc",x"cc",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"cc",x"ac",x"f0",x"ec",x"f0",x"ac",x"88",x"88",x"ac",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d5",x"b1",x"b1",x"b1",x"ad",x"d1",x"fa",x"fa",x"f6",x"fe",x"fa",x"fa",x"ff",x"fa",x"fa",x"fa",x"fa",x"d5",x"d5",x"fa",x"d6",x"ad",x"64",x"84",x"88",x"88",x"a8",x"a8",x"d5",x"fe",x"d5",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"ad",x"ad",x"b1",x"b1",x"d1",x"d1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"fd",x"fd",x"fd",x"fd",x"fe",x"d9",x"49",x"49",x"49",x"4d",x"4d",x"6d",x"6d",x"4d",x"49",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"4d",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"4d",x"49",x"49",x"4d",x"49",x"49",x"49",x"49",x"b1",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"ba",x"9a",x"76",x"56",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"31",x"51",x"51",x"51",x"55",x"75",x"55",x"51",x"51",x"2d",x"31",x"51",x"55",x"55",x"51",x"51",x"55",x"55",x"75",x"75",x"51",x"2d",x"31",x"2d",x"51",x"71",x"95",x"b9",x"b9",x"95",x"75",x"75",x"75",x"95",x"95",x"95",x"95",x"b6",x"b5",x"b5",x"b6",x"d6",x"f6",x"f6",x"ee",x"ca",x"c6",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"ca",x"ee",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ca",x"ca",x"ea",x"ea",x"ea",x"ee",x"ee",x"ee",x"ee",x"f2",x"ce",x"ca",x"ca",x"ca",x"c9",x"c6",x"ca",x"ee",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ea",x"ea",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"c5",x"ea",x"f6",x"fa",x"fa",x"b6",x"71",x"50",x"75",x"75",x"50",x"50",x"74",x"98",x"b9",x"96",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"6d",x"48",x"48",x"48",x"48",x"48",x"6d",x"6d",x"91",x"91",x"8d",x"8d",x"8d",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"48",x"48",x"48",x"48",x"6d",x"6d",x"6d",x"6d",x"6d",x"4c",x"48",x"48",x"48",x"31",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"ac",x"84",x"84",x"84",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"b1",x"b5",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"55",x"51",x"51",x"51",x"51",x"75",x"99",x"99",x"99",x"99",x"99",x"75",x"51",x"51",x"75",x"75",x"75",x"51",x"51",x"51",x"75",x"99",x"79",x"99",x"99",x"99",x"79",x"79",x"79",x"95",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a8",x"ac",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"a8",x"88",x"ac",x"cc",x"ec",x"cc",x"ec",x"ec",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"f0",x"f0",x"ec",x"cc",x"cc",x"ac",x"cc",x"cc",x"f0",x"f0",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"cc",x"ec",x"f0",x"d0",x"ac",x"88",x"ac",x"d0",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d5",x"d1",x"b1",x"b1",x"ad",x"d5",x"fa",x"fa",x"d5",x"fa",x"f6",x"da",x"fe",x"fa",x"f6",x"fa",x"fa",x"d5",x"d1",x"d1",x"fa",x"d6",x"88",x"84",x"88",x"88",x"a8",x"a8",x"d1",x"fe",x"fa",x"d1",x"d1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"d1",x"d1",x"d5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"fd",x"fd",x"fd",x"fd",x"fe",x"b5",x"29",x"49",x"49",x"49",x"49",x"4d",x"4d",x"49",x"29",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"4d",x"49",x"49",x"4d",x"49",x"49",x"49",x"49",x"6d",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"9a",x"76",x"32",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"31",x"51",x"51",x"51",x"31",x"31",x"31",x"2d",x"2d",x"2d",x"51",x"51",x"55",x"51",x"71",x"51",x"55",x"51",x"75",x"75",x"51",x"31",x"31",x"31",x"71",x"b6",x"f6",x"f6",x"f6",x"d6",x"b6",x"b6",x"b5",x"b6",x"d6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"ee",x"ca",x"ca",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"ca",x"ea",x"ee",x"ee",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ca",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"ee",x"ca",x"ca",x"ca",x"c9",x"c9",x"ee",x"f6",x"f6",x"f2",x"f2",x"ee",x"ee",x"ea",x"ee",x"ee",x"f6",x"f6",x"ee",x"ea",x"f6",x"f2",x"ee",x"ee",x"f2",x"f6",x"f6",x"f2",x"c9",x"ea",x"f2",x"f6",x"f6",x"d6",x"95",x"74",x"74",x"54",x"50",x"74",x"98",x"b8",x"b5",x"92",x"b2",x"b6",x"b6",x"92",x"92",x"92",x"8d",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"6d",x"68",x"48",x"48",x"48",x"48",x"6d",x"6d",x"8d",x"91",x"8d",x"8d",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"48",x"48",x"48",x"48",x"48",x"6d",x"6d",x"6d",x"6d",x"48",x"48",x"44",x"48",x"2d",x"2d",x"2d",x"2d",x"2d",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"d1",x"a8",x"80",x"84",x"84",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"ac",x"b5",x"a8",x"a0",x"a4",x"ad",x"95",x"79",x"99",x"99",x"b9",x"b9",x"b9",x"99",x"99",x"99",x"99",x"99",x"99",x"95",x"55",x"51",x"51",x"51",x"31",x"31",x"55",x"79",x"99",x"99",x"99",x"99",x"75",x"51",x"2d",x"51",x"51",x"75",x"75",x"99",x"79",x"75",x"75",x"99",x"99",x"99",x"99",x"75",x"55",x"75",x"99",x"95",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c8",x"a4",x"a8",x"ac",x"ac",x"ac",x"cc",x"ac",x"ac",x"ac",x"a8",x"88",x"a8",x"a8",x"cc",x"cc",x"cc",x"ec",x"f0",x"f0",x"ec",x"ec",x"cc",x"cc",x"ec",x"ec",x"ec",x"cc",x"cc",x"f0",x"ec",x"cc",x"ac",x"a8",x"a8",x"a8",x"ac",x"cc",x"f0",x"f0",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"ac",x"cc",x"cc",x"ec",x"f0",x"d0",x"cc",x"d0",x"f9",x"f1",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d1",x"b1",x"b1",x"ad",x"d6",x"fa",x"d6",x"f6",x"fa",x"d5",x"d6",x"fa",x"fa",x"f6",x"fa",x"f5",x"d1",x"b1",x"b1",x"d1",x"fa",x"fa",x"ad",x"64",x"88",x"88",x"88",x"d1",x"fe",x"fa",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"fe",x"fe",x"fd",x"fe",x"fe",x"fe",x"b5",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"29",x"29",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"4d",x"49",x"4d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"4d",x"6d",x"4d",x"49",x"49",x"49",x"49",x"49",x"29",x"6d",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"96",x"76",x"52",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"11",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"2d",x"51",x"51",x"72",x"76",x"95",x"71",x"51",x"51",x"51",x"31",x"2d",x"2d",x"2d",x"2d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"71",x"51",x"51",x"55",x"75",x"75",x"51",x"75",x"f6",x"f2",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"f2",x"f6",x"fa",x"f6",x"ca",x"ca",x"c9",x"ca",x"ea",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ca",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"ca",x"ca",x"ca",x"c9",x"ca",x"f6",x"f2",x"ee",x"ea",x"ea",x"ea",x"ea",x"c9",x"ea",x"ea",x"ea",x"f2",x"f2",x"ee",x"f2",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"f2",x"f6",x"ea",x"ee",x"ee",x"ee",x"f2",x"f2",x"f6",x"b5",x"95",x"98",x"b8",x"b9",x"b5",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"8d",x"8d",x"8d",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"6d",x"48",x"48",x"48",x"48",x"48",x"68",x"6d",x"8d",x"91",x"91",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"6d",x"6d",x"4c",x"48",x"48",x"48",x"48",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"31",x"31",x"31",x"31",x"31",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"d1",x"a8",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"a4",x"b1",x"b5",x"b9",x"b1",x"a8",x"8d",x"95",x"99",x"99",x"99",x"99",x"99",x"99",x"b9",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"31",x"31",x"31",x"31",x"31",x"2d",x"51",x"99",x"99",x"75",x"99",x"99",x"99",x"55",x"31",x"2d",x"2d",x"51",x"51",x"71",x"51",x"51",x"75",x"99",x"99",x"99",x"b9",x"75",x"55",x"55",x"75",x"75",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"c8",x"cc",x"cc",x"ec",x"cc",x"ac",x"ac",x"ac",x"cc",x"a8",x"a8",x"a8",x"88",x"88",x"a8",x"cc",x"cc",x"cc",x"f0",x"f0",x"f0",x"d0",x"ec",x"f0",x"cc",x"cc",x"ec",x"ec",x"cc",x"cc",x"ec",x"f0",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"f0",x"ec",x"cc",x"cc",x"cc",x"cc",x"ec",x"cc",x"cc",x"cc",x"a8",x"a8",x"ac",x"cc",x"cc",x"cc",x"cc",x"ac",x"cc",x"f5",x"f0",x"f0",x"f5",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d5",x"d5",x"d5",x"b1",x"f6",x"fa",x"d5",x"fa",x"f6",x"d5",x"d6",x"fa",x"fa",x"f6",x"fa",x"d5",x"d1",x"b1",x"ad",x"b1",x"f5",x"fa",x"d5",x"b1",x"a8",x"88",x"88",x"d5",x"fe",x"fa",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"fe",x"fe",x"fd",x"fe",x"fe",x"fe",x"fd",x"b5",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"29",x"29",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"4d",x"4d",x"6d",x"4d",x"49",x"4d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"49",x"d5",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"ba",x"9a",x"9a",x"76",x"76",x"56",x"32",x"32",x"12",x"0e",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"31",x"31",x"51",x"51",x"52",x"72",x"76",x"76",x"96",x"96",x"96",x"96",x"96",x"ba",x"ba",x"ba",x"da",x"da",x"da",x"75",x"51",x"51",x"51",x"51",x"31",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"75",x"75",x"75",x"da",x"f2",x"ee",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"ee",x"ea",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ee",x"f2",x"f6",x"f2",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ca",x"ca",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"ee",x"ee",x"ca",x"ca",x"c6",x"ca",x"f2",x"f6",x"ee",x"ea",x"ea",x"ea",x"ea",x"c9",x"ee",x"ee",x"ea",x"ca",x"ee",x"f2",x"f2",x"f2",x"c5",x"e9",x"ea",x"ea",x"ea",x"ea",x"ee",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"d5",x"d9",x"b9",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6e",x"8e",x"8d",x"6d",x"6d",x"8d",x"8d",x"8d",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"6d",x"48",x"48",x"48",x"48",x"48",x"48",x"6c",x"6d",x"6d",x"8d",x"91",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"6d",x"6d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"6d",x"6c",x"48",x"48",x"48",x"48",x"48",x"49",x"09",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f5",x"cd",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"a8",x"b9",x"9d",x"9d",x"b5",x"95",x"79",x"79",x"79",x"99",x"99",x"75",x"75",x"75",x"99",x"b9",x"99",x"79",x"99",x"99",x"99",x"75",x"31",x"31",x"31",x"31",x"2d",x"2d",x"55",x"99",x"75",x"55",x"79",x"99",x"99",x"75",x"51",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"51",x"75",x"99",x"b9",x"b9",x"b9",x"95",x"75",x"55",x"55",x"75",x"8d",x"a4",x"a4",x"a4",x"a4",x"a8",x"ec",x"f0",x"f0",x"f0",x"f0",x"ac",x"ac",x"cc",x"ec",x"ac",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"cc",x"cc",x"f0",x"f0",x"cc",x"cc",x"cc",x"f1",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"cc",x"a8",x"88",x"88",x"88",x"a8",x"88",x"88",x"cc",x"f0",x"cc",x"cc",x"cc",x"cc",x"ec",x"f0",x"f0",x"ec",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"d0",x"ec",x"ec",x"ec",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"d5",x"f5",x"f6",x"d5",x"fa",x"d5",x"d5",x"d6",x"fa",x"f6",x"f6",x"f6",x"d1",x"d1",x"b1",x"ad",x"b1",x"d1",x"d1",x"fa",x"fa",x"d1",x"ac",x"ad",x"f5",x"fa",x"fa",x"f5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"fd",x"fe",x"fe",x"fd",x"fe",x"fe",x"fe",x"f9",x"91",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"29",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"4d",x"4d",x"4d",x"6d",x"4d",x"49",x"4d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"49",x"b1",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"96",x"76",x"56",x"32",x"32",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"0e",x"12",x"12",x"0e",x"0e",x"0e",x"0d",x"0e",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"0e",x"2d",x"2d",x"2d",x"2e",x"2d",x"31",x"51",x"52",x"76",x"96",x"96",x"ba",x"da",x"da",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"75",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"51",x"75",x"fa",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"ce",x"f2",x"f2",x"f2",x"f6",x"f6",x"f2",x"ee",x"ca",x"c5",x"ca",x"f2",x"f6",x"f2",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c9",x"ca",x"ca",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ca",x"ca",x"ea",x"ea",x"ca",x"ca",x"c9",x"ee",x"ca",x"c9",x"c9",x"c5",x"ca",x"f6",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"c9",x"f2",x"f2",x"ee",x"c9",x"c5",x"f2",x"f6",x"f2",x"c5",x"c9",x"c9",x"ea",x"ea",x"ea",x"ea",x"ee",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"f6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"48",x"6d",x"6d",x"8d",x"8d",x"8d",x"91",x"91",x"8d",x"91",x"91",x"91",x"6d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"6d",x"6d",x"8d",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"48",x"48",x"48",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"6d",x"48",x"48",x"48",x"48",x"48",x"6c",x"6d",x"29",x"09",x"09",x"0d",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"84",x"80",x"84",x"84",x"80",x"a8",x"95",x"99",x"99",x"99",x"79",x"75",x"79",x"79",x"99",x"99",x"75",x"51",x"51",x"51",x"75",x"b9",x"75",x"75",x"99",x"79",x"99",x"75",x"31",x"2d",x"2d",x"2d",x"2d",x"51",x"75",x"99",x"55",x"51",x"75",x"99",x"99",x"79",x"75",x"51",x"51",x"2d",x"2d",x"31",x"51",x"75",x"99",x"b9",x"b9",x"99",x"99",x"b9",x"b9",x"75",x"55",x"55",x"71",x"a4",x"a4",x"a4",x"a4",x"cc",x"cc",x"ac",x"cc",x"f0",x"f0",x"cc",x"a8",x"cc",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"f0",x"ac",x"a8",x"a8",x"a8",x"f0",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"f1",x"a8",x"88",x"88",x"a8",x"88",x"a8",x"a8",x"cc",x"f0",x"cc",x"cc",x"cc",x"cc",x"f1",x"f0",x"f0",x"f0",x"f0",x"cc",x"a8",x"a8",x"ac",x"a8",x"a8",x"a8",x"ac",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"f5",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d1",x"f6",x"d5",x"d5",x"d6",x"f6",x"f5",x"f6",x"f6",x"d1",x"d1",x"d1",x"ad",x"b1",x"d1",x"d1",x"d5",x"f6",x"fa",x"f6",x"f5",x"f6",x"fa",x"fa",x"fa",x"d1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fe",x"fe",x"f9",x"8d",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"49",x"29",x"49",x"49",x"49",x"6d",x"6d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b1",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"de",x"da",x"ba",x"9a",x"96",x"76",x"52",x"32",x"12",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0e",x"0e",x"0e",x"0e",x"0e",x"0e",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"31",x"32",x"52",x"56",x"76",x"76",x"96",x"96",x"b6",x"da",x"da",x"de",x"de",x"de",x"de",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"71",x"2d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"4d",x"2d",x"31",x"91",x"f6",x"ea",x"ea",x"ca",x"ea",x"ea",x"ea",x"ee",x"f2",x"f2",x"f6",x"f6",x"f6",x"f2",x"f2",x"ee",x"f2",x"f2",x"f2",x"f6",x"f2",x"c9",x"c9",x"c9",x"f2",x"f2",x"ee",x"ea",x"ca",x"ca",x"ca",x"c9",x"c9",x"c5",x"c6",x"c6",x"ca",x"ea",x"ea",x"ca",x"ea",x"ea",x"ee",x"ee",x"ee",x"ca",x"ca",x"c6",x"c6",x"ca",x"ca",x"ee",x"ee",x"ca",x"c9",x"c6",x"c6",x"ce",x"f6",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"c9",x"f6",x"ea",x"ee",x"c5",x"ea",x"ee",x"f2",x"f2",x"ee",x"f2",x"ee",x"c9",x"c9",x"ea",x"ea",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ee",x"ee",x"ee",x"f2",x"d6",x"b6",x"92",x"92",x"92",x"92",x"72",x"6d",x"6d",x"69",x"48",x"48",x"6d",x"6d",x"91",x"8d",x"6d",x"8d",x"8d",x"8d",x"8d",x"8d",x"6d",x"6d",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"6d",x"6d",x"6d",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"48",x"48",x"48",x"48",x"68",x"6c",x"6d",x"6d",x"6d",x"6d",x"6d",x"48",x"48",x"28",x"48",x"ad",x"d1",x"d1",x"91",x"4d",x"09",x"09",x"09",x"09",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"cc",x"a8",x"84",x"80",x"84",x"8c",x"99",x"99",x"79",x"75",x"79",x"79",x"79",x"79",x"99",x"75",x"51",x"31",x"2d",x"31",x"75",x"99",x"55",x"75",x"79",x"79",x"99",x"79",x"55",x"51",x"51",x"51",x"51",x"75",x"95",x"75",x"51",x"51",x"75",x"79",x"99",x"99",x"79",x"75",x"75",x"51",x"51",x"51",x"55",x"75",x"99",x"b9",x"99",x"75",x"79",x"99",x"99",x"99",x"75",x"51",x"88",x"a4",x"a4",x"a4",x"c8",x"cc",x"ac",x"88",x"cc",x"f0",x"f0",x"cc",x"a8",x"cc",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"cc",x"a8",x"88",x"88",x"a8",x"d0",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"cc",x"f1",x"ac",x"a8",x"88",x"88",x"88",x"88",x"a8",x"d0",x"f0",x"cc",x"cc",x"cc",x"cc",x"f1",x"cc",x"cc",x"cc",x"d0",x"f0",x"cc",x"ac",x"ac",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f5",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d1",x"d5",x"d1",x"d5",x"d5",x"d5",x"d5",x"d5",x"d6",x"b1",x"d1",x"d1",x"ad",x"ad",x"b1",x"ad",x"d1",x"f6",x"fa",x"fa",x"f6",x"f6",x"fa",x"fa",x"fa",x"f5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fe",x"fd",x"fe",x"fe",x"d5",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"49",x"29",x"49",x"49",x"49",x"6d",x"6d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"d5",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"de",x"da",x"ba",x"9a",x"9a",x"76",x"76",x"76",x"76",x"76",x"76",x"56",x"56",x"56",x"56",x"56",x"56",x"56",x"56",x"52",x"52",x"52",x"56",x"56",x"56",x"56",x"56",x"52",x"56",x"76",x"76",x"76",x"76",x"76",x"76",x"76",x"76",x"76",x"96",x"96",x"9a",x"ba",x"ba",x"ba",x"da",x"de",x"de",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"71",x"2d",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"2d",x"31",x"b1",x"f2",x"ea",x"c9",x"c9",x"ca",x"ee",x"f2",x"f2",x"f6",x"f6",x"f6",x"f2",x"f2",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"c9",x"c9",x"c6",x"ee",x"f2",x"ee",x"ea",x"ea",x"ca",x"c6",x"c5",x"c9",x"ca",x"ca",x"ca",x"ce",x"ee",x"ce",x"ea",x"ea",x"ca",x"ea",x"ea",x"ea",x"ca",x"ca",x"ca",x"ca",x"ea",x"ce",x"ce",x"ca",x"ca",x"c6",x"c6",x"ca",x"ce",x"f2",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ca",x"f6",x"ee",x"ee",x"c9",x"ee",x"f2",x"ee",x"f2",x"f2",x"f6",x"ee",x"c9",x"c9",x"c9",x"ee",x"f2",x"ea",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ee",x"f2",x"b2",x"92",x"92",x"92",x"92",x"6e",x"6d",x"69",x"68",x"48",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6c",x"6c",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"48",x"44",x"48",x"8c",x"d1",x"f5",x"f5",x"d1",x"b1",x"91",x"4d",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"0d",x"0d",x"2d",x"0d",x"2d",x"0d",x"0d",x"0d",x"0d",x"0d",x"0d",x"09",x"09"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"d1",x"a8",x"84",x"88",x"91",x"79",x"75",x"75",x"75",x"79",x"79",x"75",x"79",x"99",x"75",x"31",x"2d",x"31",x"51",x"75",x"75",x"55",x"75",x"79",x"79",x"75",x"99",x"79",x"75",x"75",x"75",x"99",x"99",x"75",x"51",x"31",x"51",x"75",x"79",x"99",x"99",x"99",x"79",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"99",x"75",x"55",x"55",x"55",x"75",x"99",x"99",x"71",x"a4",x"a4",x"a4",x"a4",x"cc",x"cc",x"88",x"ac",x"f0",x"f0",x"ec",x"ac",x"88",x"ac",x"ec",x"cc",x"cc",x"f0",x"ec",x"cc",x"cc",x"cc",x"cc",x"ec",x"cc",x"a8",x"88",x"88",x"ac",x"d0",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"ac",x"d0",x"d0",x"cc",x"a8",x"88",x"88",x"a8",x"ac",x"d0",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"a8",x"a8",x"a8",x"ac",x"f0",x"f0",x"cc",x"ac",x"ac",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f1",x"f9",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"b1",x"d5",x"d1",x"d5",x"d1",x"d5",x"d5",x"d5",x"d5",x"b1",x"d1",x"d5",x"b1",x"ad",x"ad",x"ac",x"ad",x"d5",x"f6",x"fa",x"d6",x"d5",x"f6",x"fa",x"fa",x"f6",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"fd",x"fe",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"b5",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"49",x"29",x"49",x"49",x"49",x"6d",x"6d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"8d",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"da",x"da",x"da",x"de",x"de",x"da",x"da",x"da",x"da",x"da",x"da",x"da",x"de",x"da",x"da",x"da",x"da",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"95",x"09",x"2d",x"2d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"51",x"f6",x"ee",x"e9",x"c9",x"c9",x"ee",x"f6",x"f6",x"f6",x"f6",x"f6",x"f2",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"c5",x"ee",x"f2",x"ca",x"c9",x"ea",x"c6",x"f2",x"ee",x"ea",x"ea",x"ca",x"ca",x"c6",x"ca",x"ce",x"ee",x"f2",x"f2",x"f2",x"f2",x"ee",x"ee",x"ea",x"ea",x"ea",x"ca",x"ca",x"ca",x"ee",x"ee",x"ee",x"ca",x"ca",x"c6",x"ca",x"c6",x"c6",x"ca",x"ee",x"f2",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ca",x"f2",x"f2",x"ee",x"ee",x"f2",x"ee",x"c9",x"ce",x"f2",x"f2",x"ea",x"ca",x"c5",x"c9",x"ee",x"f2",x"c5",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"f2",x"b2",x"72",x"92",x"92",x"72",x"6e",x"6d",x"69",x"68",x"68",x"68",x"68",x"48",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"48",x"48",x"68",x"6c",x"6c",x"48",x"48",x"48",x"48",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"48",x"44",x"68",x"d1",x"f5",x"d1",x"d1",x"f1",x"f5",x"f9",x"d5",x"91",x"4d",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"cd",x"ad",x"71",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"95",x"71",x"71",x"75",x"79",x"75",x"55",x"51",x"75",x"79",x"79",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"31",x"51",x"55",x"79",x"79",x"79",x"75",x"79",x"79",x"79",x"75",x"79",x"99",x"75",x"55",x"79",x"99",x"51",x"31",x"51",x"51",x"55",x"75",x"99",x"75",x"8c",x"a4",x"a4",x"c8",x"cc",x"a8",x"88",x"d0",x"ec",x"ec",x"cc",x"a8",x"88",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"cc",x"cc",x"cc",x"ec",x"f0",x"d0",x"cc",x"cc",x"d0",x"cc",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"cc",x"cc",x"d0",x"d0",x"d0",x"d0",x"d0",x"d0",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"f0",x"ac",x"88",x"88",x"88",x"cc",x"f0",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"f0",x"f0",x"ec",x"ec",x"cc",x"cc",x"cc",x"cc",x"d1",x"f5",x"f9",x"fd",x"fd",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"d5",x"b1",x"b1",x"d5",x"d1",x"d5",x"d1",x"d5",x"d5",x"d5",x"d5",x"ad",x"ad",x"d1",x"b1",x"ad",x"ad",x"ad",x"ad",x"b1",x"d1",x"f6",x"f6",x"d5",x"f6",x"fa",x"f6",x"fa",x"fa",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fe",x"fd",x"fd",x"fe",x"fe",x"fe",x"fa",x"f9",x"b1",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"29",x"29",x"49",x"49",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"91",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"09",x"09",x"2d",x"2d",x"2d",x"2d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"71",x"f6",x"ea",x"ea",x"c9",x"ca",x"f2",x"f6",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ca",x"c9",x"c9",x"c5",x"ce",x"f2",x"ca",x"c9",x"c9",x"c5",x"f2",x"f2",x"ca",x"ca",x"ca",x"ce",x"f2",x"f6",x"f6",x"f6",x"f2",x"f2",x"f2",x"f2",x"f6",x"f6",x"f2",x"ee",x"ea",x"ee",x"ee",x"ee",x"ea",x"ca",x"ca",x"c9",x"c5",x"c6",x"c6",x"ca",x"ce",x"f2",x"f2",x"f2",x"e9",x"ee",x"ee",x"ea",x"ea",x"ea",x"c9",x"ee",x"f2",x"f2",x"f2",x"ee",x"ea",x"c5",x"c9",x"ee",x"ee",x"ea",x"ca",x"c5",x"c9",x"ee",x"ee",x"c5",x"ea",x"ee",x"ee",x"ea",x"ea",x"ea",x"c9",x"c5",x"ea",x"f2",x"b2",x"72",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"68",x"68",x"48",x"48",x"48",x"48",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"48",x"48",x"48",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6c",x"48",x"48",x"48",x"48",x"48",x"24",x"6c",x"d5",x"f5",x"d1",x"d1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"b1",x"91",x"6d",x"4d",x"2d",x"29",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"2d",x"2d"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"d1",x"95",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"51",x"75",x"79",x"79",x"75",x"51",x"51",x"75",x"75",x"55",x"51",x"31",x"31",x"31",x"51",x"75",x"99",x"99",x"99",x"99",x"99",x"79",x"79",x"79",x"99",x"99",x"75",x"55",x"75",x"99",x"55",x"2d",x"31",x"31",x"51",x"75",x"95",x"99",x"71",x"a4",x"a0",x"a8",x"cc",x"ac",x"ac",x"d0",x"ec",x"cc",x"ac",x"88",x"a8",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"a8",x"a8",x"ac",x"cc",x"d0",x"d0",x"d0",x"d0",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"cc",x"cc",x"ac",x"ac",x"a8",x"cc",x"f0",x"cc",x"cc",x"cc",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"cc",x"c8",x"c8",x"cc",x"cc",x"f1",x"f5",x"f9",x"f9",x"fd",x"f9",x"d5",x"f5",x"f5",x"f5",x"d5",x"ad",x"ad",x"d1",x"b1",x"d1",x"d1",x"d5",x"d1",x"d1",x"d5",x"ad",x"ad",x"b1",x"b1",x"ad",x"ad",x"ad",x"ad",x"ad",x"b1",x"d1",x"d1",x"d1",x"d5",x"f6",x"f6",x"f6",x"fa",x"fe",x"fe",x"fe",x"fd",x"f9",x"fa",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"f9",x"f9",x"91",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"29",x"29",x"49",x"49",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"49",x"8d",x"d5",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"91",x"2d",x"09",x"0d",x"2d",x"2d",x"2d",x"2d",x"31",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"51",x"91",x"f2",x"ea",x"ea",x"c6",x"ee",x"f2",x"f2",x"ea",x"ea",x"ea",x"ee",x"ee",x"ee",x"f2",x"f2",x"ee",x"c9",x"c9",x"c5",x"ca",x"f2",x"f2",x"c5",x"c9",x"c9",x"c5",x"f2",x"f2",x"ca",x"ca",x"ee",x"f2",x"f6",x"f6",x"f2",x"f2",x"f2",x"ee",x"ee",x"ee",x"f2",x"f2",x"f6",x"f2",x"ee",x"ea",x"ea",x"ea",x"ca",x"c6",x"ca",x"c9",x"c9",x"c6",x"ca",x"ce",x"ee",x"ee",x"ee",x"f2",x"e9",x"ea",x"ea",x"ea",x"ea",x"ea",x"c9",x"ca",x"ee",x"ee",x"ee",x"ee",x"ea",x"c5",x"c9",x"ee",x"ee",x"ca",x"c9",x"c5",x"c9",x"ee",x"f2",x"c6",x"ea",x"ee",x"ee",x"ea",x"ea",x"c6",x"c5",x"c5",x"ee",x"d2",x"8d",x"6d",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"48",x"48",x"48",x"48",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6c",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"6c",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"28",x"68",x"d5",x"f5",x"d5",x"d1",x"d1",x"d5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"d5",x"d1",x"b1",x"91",x"91",x"91",x"71",x"71",x"71",x"71",x"71",x"71",x"71",x"91",x"91",x"91"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"b5",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"51",x"55",x"55",x"51",x"51",x"51",x"51",x"51",x"75",x"79",x"79",x"75",x"51",x"2d",x"51",x"51",x"2d",x"2d",x"2d",x"31",x"31",x"51",x"99",x"b9",x"b9",x"b9",x"b9",x"99",x"79",x"75",x"79",x"79",x"79",x"55",x"51",x"75",x"99",x"95",x"51",x"31",x"2d",x"31",x"51",x"75",x"99",x"55",x"88",x"84",x"a8",x"cc",x"d0",x"d0",x"cc",x"cc",x"cc",x"a8",x"88",x"a8",x"cc",x"f0",x"cc",x"cc",x"cc",x"f0",x"f0",x"cc",x"ac",x"cc",x"cc",x"a8",x"ac",x"ac",x"ac",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"a8",x"a8",x"ac",x"cc",x"cc",x"cc",x"ac",x"cc",x"cc",x"d0",x"cc",x"cc",x"cc",x"d0",x"cc",x"cc",x"cc",x"cc",x"f0",x"f0",x"cc",x"ac",x"cc",x"ec",x"f0",x"ec",x"cc",x"cc",x"cc",x"cc",x"c8",x"cc",x"d0",x"f9",x"fd",x"f9",x"f5",x"f5",x"f5",x"f5",x"d5",x"b1",x"ad",x"b1",x"b1",x"b1",x"d1",x"d1",x"b1",x"b1",x"d5",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"d1",x"d1",x"ac",x"ad",x"ad",x"ad",x"ad",x"b1",x"d5",x"fa",x"f5",x"f6",x"f9",x"fe",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fe",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"f5",x"f9",x"91",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"29",x"29",x"49",x"49",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"8d",x"f6",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"71",x"2d",x"09",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"31",x"31",x"51",x"2d",x"71",x"f6",x"ee",x"ea",x"ea",x"ca",x"f2",x"f2",x"ee",x"ea",x"ea",x"ea",x"ee",x"ea",x"ee",x"f2",x"f6",x"f2",x"c9",x"c9",x"c9",x"ee",x"f2",x"ee",x"c5",x"c9",x"ca",x"c5",x"f2",x"f2",x"c9",x"ce",x"f6",x"f6",x"f2",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"f2",x"f6",x"ee",x"c6",x"c6",x"c6",x"ca",x"ca",x"ca",x"ea",x"ca",x"ca",x"f2",x"f2",x"ee",x"ea",x"ca",x"f2",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"ee",x"ee",x"ee",x"ee",x"ca",x"c6",x"ca",x"ee",x"ee",x"c9",x"c9",x"c5",x"c9",x"cd",x"f2",x"c6",x"ea",x"ee",x"ea",x"ea",x"ea",x"c5",x"c9",x"ca",x"f2",x"b1",x"6d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b1",x"8d",x"6d",x"6d",x"6d",x"48",x"48",x"48",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"d5",x"f5",x"f5",x"f5",x"d1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"b5",x"75",x"55",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"51",x"31",x"51",x"31",x"31",x"51",x"75",x"75",x"75",x"75",x"75",x"55",x"51",x"31",x"31",x"31",x"2d",x"31",x"31",x"55",x"75",x"b9",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"75",x"79",x"79",x"75",x"51",x"55",x"75",x"79",x"75",x"51",x"2d",x"2d",x"31",x"75",x"99",x"55",x"6d",x"84",x"a4",x"ac",x"cc",x"cc",x"ac",x"a8",x"a8",x"88",x"88",x"cc",x"f0",x"cc",x"cc",x"ac",x"a8",x"cc",x"f0",x"cc",x"a8",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"d0",x"ac",x"a8",x"a8",x"a8",x"cc",x"f0",x"cc",x"cc",x"cc",x"cc",x"c8",x"cc",x"a8",x"ac",x"d5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"ad",x"8d",x"8d",x"ad",x"ad",x"b1",x"ad",x"ad",x"b1",x"ad",x"8d",x"8c",x"ad",x"d1",x"f5",x"f5",x"f5",x"d5",x"d5",x"d1",x"b1",x"ad",x"ad",x"ad",x"d1",x"fa",x"f6",x"f5",x"f9",x"fe",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fd",x"f9",x"f5",x"f9",x"8d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"29",x"49",x"49",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"49",x"b1",x"d6",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ba",x"71",x"09",x"09",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"91",x"f2",x"ee",x"ea",x"ea",x"ca",x"f2",x"f2",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"f2",x"f2",x"c9",x"ca",x"ca",x"ca",x"ee",x"f2",x"f2",x"ee",x"ce",x"ee",x"ee",x"ee",x"f2",x"ee",x"c6",x"ee",x"f6",x"ee",x"ea",x"ea",x"ea",x"e9",x"ca",x"c9",x"ca",x"c5",x"ea",x"ea",x"ee",x"f2",x"f6",x"c5",x"a6",x"ca",x"ea",x"ca",x"ea",x"ea",x"ca",x"ca",x"ee",x"ee",x"f2",x"f2",x"f2",x"f6",x"f2",x"ee",x"ea",x"ca",x"c9",x"c9",x"c6",x"c9",x"ea",x"ee",x"ee",x"ea",x"ca",x"c5",x"c9",x"ea",x"ee",x"c9",x"c5",x"c5",x"ca",x"f2",x"ee",x"c5",x"ea",x"ea",x"ea",x"ea",x"ea",x"ed",x"f2",x"ee",x"ce",x"8d",x"4d",x"4d",x"4d",x"6d",x"8d",x"b1",x"d5",x"f5",x"ad",x"49",x"6d",x"6d",x"6d",x"6d",x"68",x"48",x"48",x"48",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"24",x"48",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"95",x"55",x"75",x"75",x"99",x"99",x"99",x"75",x"75",x"75",x"75",x"55",x"51",x"31",x"51",x"51",x"51",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"51",x"51",x"51",x"51",x"51",x"55",x"75",x"99",x"99",x"75",x"55",x"55",x"75",x"95",x"99",x"99",x"75",x"79",x"79",x"75",x"51",x"51",x"55",x"79",x"79",x"75",x"51",x"51",x"51",x"75",x"99",x"51",x"51",x"84",x"84",x"a8",x"ac",x"a8",x"a8",x"a8",x"88",x"88",x"a8",x"cc",x"f0",x"cc",x"ac",x"88",x"88",x"cc",x"ec",x"cc",x"a8",x"cc",x"cc",x"cc",x"ac",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"a8",x"a8",x"a8",x"88",x"a8",x"88",x"88",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"ac",x"a8",x"a8",x"a8",x"ac",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"cc",x"ac",x"88",x"88",x"88",x"ac",x"d0",x"d0",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"ac",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"b1",x"b1",x"ad",x"8d",x"ad",x"ad",x"ac",x"ad",x"ad",x"ad",x"ad",x"d1",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"d1",x"b1",x"b1",x"ad",x"b1",x"d6",x"fa",x"f6",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"f9",x"f5",x"f9",x"8d",x"25",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"28",x"49",x"49",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"48",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"4d",x"6d",x"b1",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ba",x"71",x"2d",x"0d",x"09",x"0d",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"51",x"d2",x"f2",x"ea",x"ea",x"ea",x"ea",x"f2",x"ee",x"ca",x"c9",x"ea",x"ea",x"ea",x"ea",x"f2",x"f2",x"ca",x"ca",x"ee",x"ee",x"f6",x"f6",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f6",x"ee",x"ca",x"ce",x"f6",x"e9",x"ea",x"ea",x"c9",x"c9",x"ca",x"ee",x"f2",x"ee",x"ca",x"ea",x"ea",x"f2",x"f6",x"c5",x"ce",x"ee",x"f2",x"f2",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"f2",x"f6",x"f2",x"f2",x"f6",x"ee",x"ee",x"ee",x"ea",x"ca",x"ca",x"c5",x"ca",x"ee",x"ee",x"ea",x"ca",x"c5",x"c9",x"ea",x"ee",x"c9",x"c9",x"ca",x"ee",x"f2",x"ea",x"c5",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"ee",x"ea",x"ae",x"6d",x"6d",x"8d",x"91",x"91",x"b1",x"f5",x"f5",x"f5",x"d1",x"6d",x"4d",x"6d",x"8d",x"6d",x"6d",x"6d",x"68",x"48",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"24",x"8c",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d5",x"f5",x"d5",x"f5",x"f5",x"b5",x"55",x"55",x"95",x"b9",x"b9",x"b9",x"b9",x"99",x"75",x"55",x"75",x"75",x"51",x"55",x"51",x"51",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"55",x"55",x"55",x"75",x"75",x"75",x"99",x"99",x"75",x"51",x"31",x"31",x"31",x"55",x"99",x"99",x"75",x"75",x"79",x"75",x"51",x"51",x"51",x"75",x"75",x"99",x"99",x"95",x"95",x"99",x"75",x"51",x"31",x"88",x"84",x"a4",x"a8",x"88",x"88",x"88",x"88",x"88",x"ac",x"d0",x"d0",x"a8",x"a8",x"88",x"a8",x"cc",x"cc",x"ac",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"88",x"88",x"a8",x"cc",x"d0",x"cc",x"cc",x"cc",x"cc",x"c8",x"a8",x"a8",x"88",x"ac",x"fa",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d1",x"ad",x"8d",x"8d",x"ad",x"ad",x"b1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d1",x"ad",x"b1",x"f6",x"f6",x"fa",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"f5",x"f5",x"f9",x"b1",x"25",x"24",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"28",x"49",x"49",x"49",x"4d",x"4d",x"49",x"4d",x"4d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"6d",x"d5",x"d5",x"d5",x"d5",x"b1",x"b1",x"d5",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"d9",x"4d",x"09",x"09",x"09",x"09",x"29",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"91",x"f2",x"ee",x"ee",x"ea",x"ea",x"ea",x"ee",x"ce",x"c5",x"c5",x"ca",x"ca",x"ea",x"ea",x"ee",x"f2",x"f2",x"f2",x"f6",x"f2",x"f6",x"fa",x"f6",x"f2",x"f2",x"f2",x"f2",x"f2",x"f6",x"f2",x"ce",x"ce",x"f6",x"ea",x"ea",x"c9",x"ca",x"ca",x"f2",x"fa",x"fa",x"f6",x"ca",x"c6",x"ca",x"ee",x"f2",x"c6",x"f6",x"f6",x"f6",x"fa",x"f6",x"f6",x"f6",x"f6",x"fa",x"f6",x"f2",x"ee",x"ea",x"ea",x"f6",x"ee",x"f2",x"f2",x"f2",x"ee",x"ee",x"ca",x"c5",x"ea",x"ea",x"ea",x"ca",x"c9",x"c5",x"ca",x"ea",x"c9",x"ca",x"ee",x"f2",x"ee",x"ea",x"c9",x"ea",x"ea",x"ea",x"ee",x"ee",x"ca",x"c5",x"c5",x"8d",x"71",x"b1",x"d5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"b1",x"48",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6c",x"48",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6c",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"24",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d5",x"f5",x"f5",x"75",x"55",x"75",x"99",x"99",x"75",x"75",x"95",x"99",x"75",x"55",x"75",x"75",x"75",x"75",x"75",x"55",x"75",x"75",x"95",x"99",x"b9",x"b9",x"99",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"99",x"51",x"31",x"31",x"31",x"31",x"51",x"75",x"99",x"75",x"75",x"75",x"75",x"55",x"51",x"51",x"51",x"51",x"75",x"75",x"75",x"75",x"75",x"51",x"2d",x"31",x"68",x"a4",x"a8",x"ac",x"88",x"88",x"88",x"a8",x"a8",x"cc",x"d0",x"ac",x"88",x"88",x"ac",x"cc",x"ec",x"cc",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"ac",x"ac",x"cc",x"cc",x"f0",x"f0",x"f0",x"ec",x"cc",x"cc",x"ac",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"ac",x"cc",x"cc",x"cc",x"cc",x"ac",x"ac",x"d0",x"d0",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"d1",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d5",x"d5",x"d1",x"d1",x"d5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"d1",x"ad",x"b1",x"d5",x"f9",x"f9",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fe",x"fe",x"f5",x"f5",x"f5",x"d5",x"b1",x"6d",x"49",x"24",x"24",x"25",x"25",x"25",x"29",x"29",x"28",x"29",x"29",x"29",x"49",x"49",x"6d",x"6d",x"49",x"49",x"4d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"d5",x"fa",x"fa",x"fa",x"fa",x"f6",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"b9",x"71",x"4d",x"09",x"09",x"09",x"09",x"09",x"0d",x"09",x"6d",x"d2",x"f2",x"ee",x"ea",x"ea",x"ea",x"ee",x"ce",x"ca",x"c6",x"ca",x"c9",x"c9",x"ea",x"ca",x"ca",x"ee",x"f2",x"ee",x"f2",x"f6",x"f6",x"f2",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"ca",x"f6",x"ee",x"c9",x"c9",x"ca",x"ca",x"ee",x"f2",x"ee",x"f2",x"f2",x"ca",x"ca",x"ee",x"f2",x"f2",x"f2",x"ee",x"ee",x"ee",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ee",x"ea",x"c5",x"c9",x"f6",x"f2",x"f2",x"ee",x"ee",x"ee",x"ee",x"ee",x"ce",x"ea",x"ea",x"ea",x"ca",x"c5",x"c5",x"c6",x"ea",x"ee",x"ee",x"ee",x"ee",x"ea",x"ca",x"c5",x"ea",x"ea",x"ea",x"ee",x"ca",x"c6",x"c5",x"d1",x"d5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"d1",x"d1",x"8d",x"48",x"48",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"48",x"6d",x"6d",x"6d",x"6c",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6c",x"48",x"48",x"48",x"44",x"24",x"24",x"b1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"b5",x"75",x"75",x"99",x"99",x"55",x"31",x"31",x"75",x"99",x"75",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"99",x"b9",x"b9",x"99",x"99",x"75",x"75",x"75",x"75",x"75",x"75",x"75",x"99",x"99",x"51",x"2d",x"31",x"31",x"2d",x"51",x"75",x"99",x"75",x"75",x"75",x"75",x"55",x"31",x"2d",x"51",x"31",x"31",x"51",x"51",x"51",x"51",x"31",x"2d",x"11",x"8d",x"a8",x"a8",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"d0",x"cc",x"ac",x"a8",x"ac",x"cc",x"cc",x"cc",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d1",x"ad",x"b1",x"d1",x"f5",x"fe",x"fd",x"fd",x"fd",x"fd",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fe",x"f9",x"f5",x"f5",x"f9",x"f5",x"d1",x"91",x"6d",x"49",x"49",x"49",x"49",x"29",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"4d",x"4d",x"49",x"4d",x"4d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"8d",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"da",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"b5",x"71",x"4d",x"2d",x"2d",x"2d",x"0d",x"09",x"b1",x"f2",x"ee",x"ea",x"ea",x"ea",x"ca",x"ee",x"ce",x"ca",x"c6",x"ca",x"c9",x"c9",x"ca",x"ca",x"c5",x"ca",x"ee",x"ee",x"f2",x"f6",x"f2",x"ee",x"ee",x"ea",x"ea",x"ee",x"ee",x"ea",x"ea",x"ee",x"f2",x"c9",x"f2",x"f2",x"c9",x"c9",x"c6",x"ca",x"ea",x"e9",x"c5",x"f2",x"f2",x"ca",x"ca",x"ee",x"f2",x"f6",x"ca",x"c5",x"c9",x"ea",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"ca",x"c5",x"c9",x"f6",x"f2",x"f2",x"ee",x"ee",x"ca",x"ca",x"ee",x"ee",x"ee",x"ea",x"ca",x"c5",x"c5",x"ca",x"ca",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"ca",x"c5",x"ea",x"ca",x"ee",x"ee",x"c5",x"c6",x"cd",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d1",x"f5",x"d5",x"6c",x"48",x"48",x"68",x"6c",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"6d",x"6c",x"6c",x"6c",x"6d",x"6d",x"6c",x"6d",x"8d",x"91",x"b6",x"b6",x"b6",x"91",x"91",x"6d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6c",x"68",x"48",x"48",x"48",x"44",x"48",x"8c",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"95",x"55",x"79",x"99",x"51",x"31",x"31",x"2d",x"75",x"99",x"75",x"55",x"55",x"75",x"55",x"55",x"55",x"75",x"75",x"99",x"99",x"75",x"75",x"75",x"95",x"99",x"99",x"75",x"55",x"55",x"75",x"75",x"75",x"75",x"79",x"51",x"2d",x"2d",x"2d",x"2d",x"51",x"99",x"79",x"51",x"75",x"75",x"75",x"55",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"51",x"2d",x"2d",x"0d",x"b1",x"ac",x"a8",x"a8",x"a8",x"ac",x"ac",x"ac",x"a8",x"cc",x"d0",x"d0",x"d0",x"d0",x"d1",x"cc",x"ac",x"a8",x"ac",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"f0",x"f0",x"f0",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"f0",x"d0",x"cc",x"cc",x"d0",x"f1",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"ac",x"a8",x"a8",x"ac",x"cc",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"ad",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"d5",x"ad",x"8d",x"d1",x"fe",x"fd",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fe",x"fe",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"d5",x"b1",x"8d",x"6d",x"49",x"24",x"24",x"24",x"24",x"29",x"49",x"49",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b1",x"fa",x"f6",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"d5",x"d2",x"d6",x"d6",x"d6",x"d6",x"d6",x"d1",x"b1",x"d1",x"da",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"b5",x"71",x"4d",x"4d",x"d2",x"ee",x"ea",x"ea",x"ea",x"ea",x"c9",x"ea",x"ee",x"ce",x"c5",x"c6",x"c9",x"ca",x"ca",x"ca",x"c6",x"c6",x"ca",x"f2",x"f6",x"f2",x"ee",x"ea",x"ea",x"ea",x"ea",x"ee",x"ea",x"ea",x"ea",x"ee",x"f2",x"ca",x"ee",x"f6",x"ee",x"ca",x"c5",x"c5",x"c5",x"ca",x"ca",x"f6",x"ee",x"ca",x"ca",x"ee",x"f6",x"f2",x"c5",x"c9",x"c9",x"ea",x"ee",x"ee",x"ee",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"ee",x"fa",x"f2",x"ee",x"f6",x"ee",x"c6",x"c6",x"c6",x"ce",x"f2",x"ee",x"ca",x"c5",x"c9",x"ee",x"f2",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"c6",x"ea",x"c6",x"ee",x"ee",x"c6",x"c9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"b1",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"6d",x"48",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"48",x"68",x"6c",x"6d",x"6d",x"6c",x"6c",x"48",x"48",x"48",x"48",x"28",x"24",x"48",x"ac",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"75",x"55",x"99",x"75",x"2d",x"2d",x"2d",x"51",x"75",x"75",x"55",x"51",x"55",x"55",x"55",x"55",x"55",x"75",x"99",x"99",x"75",x"51",x"51",x"51",x"55",x"75",x"99",x"79",x"75",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"71",x"51",x"55",x"75",x"75",x"75",x"51",x"51",x"75",x"75",x"55",x"51",x"51",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"51",x"31",x"2d",x"2d",x"2d",x"b1",x"ac",x"a8",x"a8",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"cc",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"f0",x"f0",x"cc",x"cc",x"d0",x"f0",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"cc",x"ac",x"ac",x"ac",x"ac",x"cc",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"a8",x"a8",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"f5",x"f9",x"f9",x"f5",x"f5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"f9",x"d5",x"d5",x"f9",x"fa",x"f9",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d5",x"d5",x"d5",x"b1",x"b1",x"91",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"24",x"29",x"91",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f5",x"f9",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"d5",x"d5",x"b1",x"b1",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d1",x"d1",x"d1",x"b1",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"da",x"d6",x"f2",x"ee",x"ea",x"ea",x"ea",x"ea",x"c9",x"c9",x"ee",x"f2",x"ee",x"ce",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ee",x"f6",x"f2",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"ea",x"ea",x"c5",x"ee",x"f2",x"ca",x"ca",x"f2",x"f2",x"f2",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"ea",x"c5",x"ca",x"f2",x"f6",x"f6",x"c9",x"c9",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"e9",x"c9",x"c9",x"f2",x"f2",x"ee",x"c9",x"f2",x"f2",x"ca",x"a5",x"c6",x"ca",x"ee",x"ee",x"ee",x"ca",x"ee",x"ee",x"ee",x"ea",x"ca",x"ca",x"ea",x"ea",x"ea",x"c6",x"c5",x"ca",x"c5",x"ee",x"ea",x"c6",x"cd",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"8d",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"48",x"6c",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6c",x"91",x"fb",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"b6",x"6d",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"24",x"24",x"48",x"8c",x"b1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"51",x"55",x"99",x"75",x"2d",x"51",x"51",x"75",x"75",x"51",x"51",x"51",x"75",x"55",x"55",x"55",x"51",x"75",x"99",x"75",x"51",x"31",x"31",x"31",x"31",x"55",x"79",x"99",x"75",x"55",x"75",x"55",x"55",x"55",x"75",x"75",x"75",x"75",x"75",x"99",x"75",x"51",x"51",x"51",x"75",x"55",x"51",x"51",x"51",x"51",x"31",x"31",x"2d",x"31",x"31",x"51",x"2d",x"2d",x"2d",x"2d",x"b1",x"ac",x"a8",x"a8",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"ac",x"a8",x"88",x"a8",x"a8",x"a8",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"f0",x"cc",x"a8",x"ac",x"ac",x"d0",x"f0",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f1",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"ec",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"88",x"a8",x"88",x"88",x"a8",x"a8",x"a8",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"84",x"d5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fa",x"f9",x"fd",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"f9",x"fa",x"f5",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"b1",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"25",x"49",x"6d",x"d5",x"fa",x"f9",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"d6",x"b1",x"b1",x"b1",x"b1",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d1",x"d1",x"d1",x"ad",x"d6",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f6",x"ee",x"ee",x"ea",x"ea",x"ea",x"ca",x"ca",x"c5",x"ea",x"f2",x"f2",x"ee",x"ee",x"ee",x"ee",x"ce",x"ea",x"ee",x"f2",x"f6",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"c5",x"ee",x"f2",x"c5",x"ca",x"ee",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"c9",x"c9",x"ee",x"f2",x"f2",x"f6",x"f2",x"ea",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"e9",x"c9",x"c9",x"c9",x"ee",x"ee",x"ca",x"c9",x"f2",x"f2",x"ca",x"c5",x"ca",x"ca",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ca",x"ca",x"ca",x"ca",x"ea",x"ea",x"c5",x"c5",x"c5",x"c6",x"ea",x"ea",x"c9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"d1",x"6c",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"6d",x"6d",x"6d",x"6d",x"6d",x"68",x"8d",x"da",x"fb",x"f5",x"f5",x"f6",x"f6",x"fa",x"fa",x"fe",x"ff",x"b6",x"68",x"48",x"48",x"48",x"28",x"24",x"48",x"48",x"48",x"8c",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"51",x"55",x"75",x"99",x"75",x"95",x"95",x"75",x"51",x"51",x"51",x"51",x"51",x"55",x"55",x"55",x"51",x"75",x"75",x"51",x"31",x"31",x"31",x"31",x"2d",x"51",x"75",x"99",x"71",x"55",x"55",x"55",x"55",x"55",x"31",x"51",x"75",x"75",x"75",x"51",x"51",x"31",x"51",x"51",x"75",x"51",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"2d",x"2d",x"2d",x"2d",x"4d",x"cd",x"a8",x"88",x"a8",x"a8",x"a8",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"c8",x"cc",x"f0",x"f0",x"a8",x"a8",x"88",x"88",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f1",x"a8",x"a8",x"88",x"a8",x"a8",x"88",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"84",x"d5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"d5",x"f5",x"f5",x"f5",x"f9",x"fe",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"f5",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"d5",x"69",x"04",x"24",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"24",x"24",x"6d",x"d5",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"da",x"d6",x"f6",x"d6",x"d5",x"d5",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d1",x"b1",x"b1",x"b1",x"b1",x"d6",x"d5",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f2",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"c9",x"ca",x"ca",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f6",x"ee",x"ea",x"ea",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"c9",x"c5",x"c9",x"ee",x"ee",x"c5",x"c9",x"ee",x"ee",x"ee",x"f2",x"f2",x"ee",x"ee",x"ee",x"ea",x"c5",x"ce",x"f6",x"f2",x"ea",x"ea",x"f6",x"f2",x"ca",x"ca",x"ea",x"ee",x"ea",x"ea",x"ea",x"c9",x"c5",x"c5",x"c9",x"ea",x"ee",x"c9",x"f2",x"f6",x"ee",x"c6",x"e9",x"ee",x"ca",x"c9",x"ca",x"ee",x"ee",x"c9",x"c5",x"ee",x"ee",x"ea",x"ea",x"ea",x"ca",x"c6",x"c5",x"c5",x"c6",x"ea",x"ea",x"ed",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"6c",x"24",x"28",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"48",x"b6",x"ff",x"f5",x"f6",x"f6",x"f6",x"f6",x"fa",x"fa",x"fa",x"fa",x"ff",x"91",x"48",x"44",x"44",x"24",x"24",x"48",x"8d",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d5",x"51",x"51",x"51",x"55",x"75",x"71",x"51",x"51",x"31",x"2d",x"51",x"51",x"51",x"51",x"55",x"51",x"51",x"75",x"75",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"51",x"75",x"75",x"51",x"55",x"55",x"55",x"55",x"51",x"31",x"31",x"51",x"51",x"51",x"51",x"2d",x"31",x"51",x"51",x"51",x"51",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"2d",x"2d",x"2d",x"2d",x"0d",x"6d",x"cd",x"ac",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"a8",x"a8",x"a8",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"f0",x"cc",x"ac",x"ac",x"ac",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"88",x"88",x"88",x"88",x"88",x"a8",x"cc",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"a8",x"cc",x"cc",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"84",x"d5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"fd",x"f9",x"f9",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"f5",x"f5",x"f9",x"f5",x"f5",x"f9",x"f9",x"fa",x"f9",x"f9",x"91",x"49",x"49",x"49",x"49",x"29",x"25",x"25",x"24",x"25",x"29",x"49",x"91",x"d5",x"fa",x"f9",x"f9",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"f6",x"f6",x"f6",x"d6",x"d6",x"d6",x"d6",x"f6",x"d6",x"d6",x"d6",x"d2",x"b1",x"d1",x"b1",x"ad",x"d1",x"d5",x"ad",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f6",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"c9",x"c5",x"c6",x"ea",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"ce",x"c9",x"ee",x"ee",x"ee",x"c5",x"c9",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"c9",x"f2",x"f2",x"ee",x"c5",x"c9",x"f2",x"ee",x"ca",x"ca",x"ea",x"ee",x"ea",x"ea",x"ee",x"ee",x"ea",x"ca",x"c9",x"c9",x"ea",x"f2",x"f2",x"ee",x"ca",x"ee",x"ee",x"c9",x"c6",x"ca",x"ca",x"ca",x"ca",x"c9",x"ca",x"ca",x"ee",x"ea",x"ee",x"ee",x"ea",x"ea",x"ea",x"ca",x"ea",x"ca",x"ee",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"91",x"8c",x"68",x"48",x"44",x"24",x"24",x"24",x"24",x"48",x"48",x"48",x"48",x"24",x"8d",x"fa",x"ff",x"d1",x"d1",x"d1",x"d5",x"d5",x"d5",x"f6",x"fa",x"fa",x"fe",x"db",x"48",x"24",x"68",x"8c",x"ad",x"b1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"b5",x"51",x"51",x"31",x"31",x"51",x"2d",x"2d",x"2d",x"2d",x"2d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"55",x"75",x"51",x"2d",x"31",x"2d",x"31",x"31",x"55",x"75",x"51",x"51",x"51",x"55",x"51",x"51",x"51",x"51",x"2d",x"2d",x"2d",x"2d",x"2d",x"31",x"51",x"51",x"51",x"51",x"51",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"b1",x"d1",x"ac",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"c8",x"cc",x"c8",x"cc",x"cc",x"a8",x"cc",x"f0",x"d0",x"ac",x"ac",x"cc",x"cc",x"ac",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"ac",x"ac",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"cc",x"a8",x"a8",x"cc",x"cc",x"cc",x"a8",x"ac",x"cc",x"a8",x"c8",x"cc",x"cc",x"c8",x"c8",x"cc",x"a8",x"cc",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"f5",x"f5",x"f5",x"f5",x"f9",x"fd",x"fd",x"fe",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"fd",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"f5",x"f5",x"f9",x"f5",x"f5",x"fa",x"f5",x"f9",x"f9",x"d5",x"91",x"91",x"8d",x"6d",x"6d",x"49",x"49",x"48",x"49",x"6d",x"b1",x"f9",x"f9",x"fa",x"fa",x"f9",x"fa",x"f9",x"fa",x"f6",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"f6",x"f6",x"f6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d1",x"d1",x"d1",x"b1",x"b1",x"d1",x"d1",x"89",x"d6",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"c9",x"ca",x"ca",x"c5",x"c6",x"ca",x"ea",x"ea",x"ee",x"ea",x"ea",x"ea",x"ee",x"f2",x"ee",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ee",x"f2",x"f2",x"ee",x"ee",x"f2",x"ee",x"ca",x"c5",x"c9",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"f2",x"f2",x"c9",x"c9",x"c9",x"ee",x"ee",x"e9",x"c9",x"ea",x"ea",x"ea",x"e9",x"f2",x"f2",x"ee",x"ca",x"c9",x"ca",x"ee",x"f2",x"ee",x"c5",x"c9",x"f2",x"ee",x"a5",x"c6",x"ca",x"ee",x"ca",x"c6",x"ca",x"ee",x"c6",x"ca",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ca",x"f1",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"8d",x"6c",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"24",x"b1",x"ff",x"fb",x"cd",x"d1",x"b1",x"b1",x"d1",x"d1",x"d1",x"f6",x"fa",x"fa",x"ff",x"8d",x"68",x"ac",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"95",x"51",x"51",x"51",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"55",x"75",x"55",x"51",x"51",x"51",x"75",x"75",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"31",x"31",x"51",x"51",x"51",x"31",x"31",x"31",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"2d",x"2d",x"2d",x"2d",x"0d",x"6d",x"d1",x"d1",x"a8",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a4",x"88",x"a8",x"a8",x"c8",x"c8",x"c8",x"a8",x"c8",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"cd",x"d0",x"cc",x"ac",x"cc",x"d0",x"cc",x"a8",x"a8",x"a8",x"c8",x"a8",x"a8",x"a8",x"a8",x"cc",x"a8",x"a8",x"c8",x"cc",x"cc",x"c8",x"c8",x"c8",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"a8",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"f5",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f5",x"f9",x"fa",x"fa",x"f9",x"f9",x"fa",x"f9",x"f9",x"d5",x"d5",x"f5",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"f5",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"d5",x"d6",x"f6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d2",x"d1",x"b1",x"d1",x"d6",x"d1",x"b1",x"d1",x"b1",x"d1",x"89",x"b1",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"c5",x"ca",x"ca",x"ca",x"ca",x"ea",x"ea",x"ee",x"ce",x"ea",x"ea",x"ee",x"f2",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"f2",x"f2",x"ce",x"ea",x"ee",x"f2",x"ee",x"ca",x"c5",x"c9",x"c9",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ca",x"f2",x"f2",x"ea",x"ca",x"ca",x"ca",x"ee",x"ee",x"c9",x"c9",x"ca",x"ea",x"ea",x"ea",x"f6",x"ee",x"ca",x"c9",x"c5",x"ca",x"f2",x"ee",x"ea",x"c9",x"c5",x"ee",x"f2",x"ea",x"c9",x"ed",x"ee",x"ca",x"c6",x"c6",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c6",x"ed",x"f5",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d1",x"b1",x"b1",x"8c",x"8c",x"8c",x"68",x"6c",x"da",x"ff",x"d6",x"ac",x"ad",x"cd",x"d1",x"d1",x"d1",x"d1",x"d1",x"f6",x"fa",x"fa",x"fa",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"91",x"51",x"51",x"51",x"31",x"31",x"2d",x"2d",x"4d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"51",x"55",x"75",x"75",x"75",x"75",x"75",x"75",x"51",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"31",x"31",x"31",x"51",x"51",x"31",x"31",x"2d",x"2d",x"2d",x"2d",x"0d",x"0d",x"4d",x"d1",x"d1",x"f1",x"ac",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"d1",x"d1",x"d1",x"d1",x"ad",x"d1",x"d1",x"d1",x"d1",x"cc",x"d1",x"d1",x"d1",x"cd",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"ac",x"cc",x"cc",x"ac",x"ac",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"ac",x"a8",x"cc",x"a8",x"a8",x"a8",x"a8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"d1",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"fe",x"fe",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f6",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"b1",x"b1",x"d6",x"d5",x"d5",x"d5",x"d6",x"d6",x"d6",x"d6",x"d6",x"d1",x"d5",x"d1",x"d1",x"d1",x"d1",x"b1",x"b1",x"d1",x"d1",x"b1",x"89",x"8d",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c5",x"c9",x"c6",x"c6",x"ca",x"ca",x"ea",x"ea",x"ca",x"ea",x"c6",x"ee",x"ee",x"ea",x"ea",x"ea",x"ca",x"c5",x"ce",x"f2",x"ee",x"c9",x"ca",x"ee",x"f2",x"ee",x"ce",x"c9",x"c5",x"c9",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"c5",x"f2",x"ee",x"ca",x"ca",x"c9",x"c9",x"ea",x"ee",x"ea",x"c9",x"c9",x"ca",x"ea",x"ea",x"f6",x"ee",x"ea",x"ca",x"ca",x"ee",x"f2",x"ee",x"ea",x"c9",x"c5",x"c9",x"f2",x"ee",x"ca",x"ea",x"ea",x"c6",x"c5",x"ca",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c6",x"c6",x"f1",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d5",x"d1",x"d1",x"b1",x"d1",x"fa",x"ff",x"d6",x"d1",x"d1",x"d1",x"d1",x"d1",x"ad",x"b1",x"d1",x"f5",x"fa",x"fe",x"fe",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"71",x"31",x"51",x"51",x"51",x"31",x"31",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"2d",x"51",x"55",x"75",x"75",x"75",x"51",x"31",x"2d",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"2d",x"31",x"31",x"31",x"31",x"31",x"31",x"31",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"4d",x"b1",x"f5",x"d1",x"f5",x"cd",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"fe",x"fe",x"fa",x"fa",x"d5",x"d6",x"fe",x"fa",x"fa",x"d1",x"fa",x"fe",x"fa",x"d5",x"b1",x"a8",x"a8",x"88",x"a8",x"a8",x"c8",x"cc",x"c8",x"c8",x"a8",x"cc",x"cc",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"a8",x"a8",x"ac",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"fa",x"f5",x"f5",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"fa",x"f9",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"d6",x"d6",x"d6",x"d6",x"d5",x"d1",x"d1",x"d1",x"b1",x"ad",x"b1",x"d1",x"d1",x"d1",x"8d",x"89",x"69",x"da",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"ea",x"c5",x"c5",x"c6",x"c6",x"c6",x"c5",x"c5",x"c5",x"c5",x"c5",x"c6",x"ca",x"ea",x"ca",x"ca",x"ea",x"ca",x"ee",x"ee",x"ea",x"ea",x"ca",x"c9",x"c5",x"ee",x"ee",x"c5",x"c5",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ca",x"c6",x"ca",x"ea",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"c5",x"f2",x"ee",x"ca",x"c9",x"c9",x"c9",x"ea",x"ee",x"ea",x"ca",x"c9",x"ca",x"ea",x"e9",x"f2",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"ea",x"c9",x"ca",x"c5",x"c9",x"f2",x"ca",x"ca",x"ca",x"ca",x"c6",x"c5",x"ea",x"ee",x"c6",x"c6",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c6",x"cd",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"fa",x"fe",x"ff",x"fb",x"fa",x"f6",x"d6",x"d6",x"d1",x"d1",x"d1",x"d1",x"f9",x"fa",x"fe",x"fa",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"6d",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"2d",x"2d",x"31",x"31",x"31",x"31",x"31",x"2d",x"2d",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"31",x"31",x"4d",x"2d",x"2d",x"31",x"51",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"0d",x"4d",x"b1",x"f5",x"f1",x"d1",x"f5",x"d1",x"88",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"ac",x"fa",x"fe",x"fe",x"ff",x"fa",x"fe",x"ff",x"ff",x"fe",x"fa",x"fe",x"ff",x"ff",x"fe",x"fe",x"fa",x"d5",x"ac",x"a8",x"c8",x"ac",x"ac",x"ac",x"ac",x"cc",x"c8",x"ac",x"a8",x"cc",x"cc",x"a8",x"88",x"88",x"a8",x"a8",x"a8",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"c8",x"cc",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"84",x"88",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"fa",x"f9",x"fa",x"fa",x"f9",x"f9",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"b1",x"8d",x"ad",x"b1",x"b1",x"b1",x"b1",x"b1",x"d1",x"d6",x"d6",x"d1",x"b1",x"b1",x"b1",x"ad",x"b1",x"d1",x"d5",x"d1",x"ad",x"8d",x"89",x"69",x"da",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ee",x"c5",x"c6",x"c6",x"c5",x"c5",x"c5",x"c5",x"c5",x"c9",x"ca",x"c6",x"c6",x"c6",x"ca",x"ca",x"ea",x"ea",x"ee",x"ee",x"ea",x"ea",x"ca",x"ca",x"c6",x"ee",x"ee",x"c5",x"c6",x"f2",x"ee",x"ee",x"ee",x"ee",x"f2",x"f2",x"ca",x"c6",x"ea",x"ea",x"ee",x"ee",x"ea",x"ea",x"ca",x"c6",x"f2",x"ee",x"ca",x"c5",x"c5",x"c9",x"c6",x"ea",x"ea",x"c9",x"c9",x"c9",x"ca",x"c9",x"c9",x"ee",x"f2",x"f2",x"ee",x"ee",x"ee",x"ea",x"c9",x"ca",x"c6",x"ca",x"ee",x"ca",x"ca",x"ca",x"ca",x"ca",x"ea",x"ea",x"ca",x"c5",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c6",x"c9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"fa",x"fa",x"fa",x"fa",x"ff",x"f6",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f5",x"f5",x"6d",x"2d",x"2d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"0d",x"2d",x"6d",x"b1",x"f5",x"f5",x"f1",x"f1",x"f5",x"d1",x"ac",x"88",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"f5",x"fe",x"fe",x"ff",x"fe",x"fe",x"ff",x"ff",x"ff",x"f9",x"fe",x"ff",x"fe",x"fe",x"fe",x"fe",x"f9",x"d5",x"cd",x"c8",x"a8",x"ac",x"cc",x"ac",x"c8",x"c8",x"a8",x"a8",x"cc",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"84",x"88",x"ad",x"f5",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"da",x"b1",x"ad",x"8d",x"8d",x"8d",x"8d",x"ad",x"b1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"b1",x"b1",x"ad",x"8d",x"89",x"89",x"69",x"da",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f6",x"ee",x"ea",x"ca",x"ca",x"ca",x"c9",x"c9",x"c6",x"c6",x"ca",x"ca",x"c9",x"ca",x"ea",x"ea",x"ea",x"ea",x"ee",x"ee",x"ea",x"ea",x"c6",x"ca",x"c6",x"ee",x"ee",x"ca",x"c6",x"f2",x"ee",x"ea",x"ca",x"ea",x"ee",x"ee",x"ee",x"c6",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"ee",x"ee",x"ee",x"ee",x"ca",x"ca",x"c9",x"ea",x"ea",x"ca",x"c9",x"ca",x"c6",x"c9",x"c5",x"ee",x"ee",x"ee",x"ee",x"ee",x"ea",x"ea",x"c9",x"ca",x"c5",x"ca",x"ee",x"ea",x"ca",x"ca",x"ea",x"ea",x"ca",x"ca",x"c6",x"c5",x"c6",x"ca",x"ca",x"ca",x"ca",x"c6",x"c6",x"ed",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fa",x"fe",x"ff",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"6d",x"2d",x"2d",x"2d",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"0d",x"4d",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"cd",x"88",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"d1",x"fa",x"fa",x"ff",x"fa",x"fa",x"ff",x"ff",x"ff",x"f5",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"d1",x"cc",x"a8",x"a8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"ac",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"f9",x"f5",x"f5",x"f9",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"d5",x"ad",x"8d",x"8d",x"8d",x"8d",x"ad",x"ad",x"ad",x"d1",x"d6",x"d5",x"d5",x"d5",x"d1",x"b1",x"ad",x"8d",x"8d",x"89",x"69",x"8d",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f6",x"ee",x"ea",x"ee",x"ea",x"e9",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ee",x"ee",x"ea",x"ca",x"ca",x"ca",x"ee",x"ee",x"ca",x"c6",x"c9",x"c6",x"c9",x"ee",x"ee",x"c9",x"ce",x"ee",x"ca",x"ca",x"ca",x"ca",x"ea",x"ee",x"c5",x"ca",x"ea",x"ea",x"ea",x"ea",x"ca",x"c6",x"ca",x"c6",x"ee",x"f2",x"f2",x"ee",x"ee",x"ee",x"ea",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"c5",x"ea",x"ea",x"ee",x"ee",x"ea",x"e9",x"ca",x"ca",x"c6",x"c5",x"ca",x"f2",x"ca",x"ea",x"ea",x"ca",x"ca",x"ca",x"ca",x"c6",x"c5",x"c6",x"ca",x"ca",x"ca",x"c6",x"c6",x"c9",x"f5",x"d5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"f5",x"f1",x"f1",x"f9",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"ff",x"ff",x"fe",x"fa",x"fe",x"fe",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"b1",x"0d",x"0d",x"2d",x"2d",x"2d",x"2d",x"31",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"0d",x"2d",x"2d",x"2d",x"0c",x"0c",x"0c",x"0d",x"0d",x"0d",x"0d",x"2d",x"91",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"ac",x"84",x"88",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"ac",x"fa",x"fe",x"fa",x"fa",x"fa",x"ff",x"ff",x"fe",x"f5",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"f5",x"f5",x"d1",x"a8",x"a8",x"ac",x"a8",x"c8",x"c8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"64",x"88",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"d6",x"d1",x"ad",x"89",x"8d",x"8d",x"8d",x"ad",x"b1",x"b1",x"b1",x"b1",x"b1",x"ad",x"8d",x"8d",x"8d",x"8d",x"89",x"65",x"b1",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f2",x"ca",x"c6",x"ea",x"ea",x"ee",x"ee",x"ea",x"ee",x"ee",x"ca",x"ca",x"ea",x"ea",x"ca",x"ca",x"ca",x"ee",x"ee",x"ca",x"c5",x"ca",x"ca",x"c6",x"ca",x"ee",x"ee",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ce",x"ee",x"c9",x"c5",x"ca",x"ea",x"ea",x"ea",x"ca",x"c6",x"c5",x"c5",x"ca",x"ca",x"ce",x"ed",x"ee",x"f2",x"c9",x"c9",x"ca",x"ca",x"c9",x"ca",x"ca",x"c9",x"ca",x"ea",x"ee",x"ee",x"ea",x"ca",x"c6",x"c6",x"c5",x"c9",x"ee",x"ee",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c6",x"c5",x"c5",x"c6",x"ca",x"c6",x"c6",x"c9",x"f1",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"d1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"f9",x"fa",x"fa",x"fa",x"fe",x"ff",x"ff",x"fe",x"ff",x"ff",x"ff",x"fe",x"ff",x"ff",x"fe",x"fe",x"fa",x"f5",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f1",x"4d",x"0d",x"0d",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"31",x"31",x"31",x"51",x"51",x"31",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"31",x"31",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"51",x"71",x"71",x"71",x"71",x"51",x"51",x"4d",x"2d",x"0d",x"2d",x"4d",x"91",x"f1",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"f1",x"f5",x"f5",x"d1",x"88",x"88",x"88",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"fa",x"fe",x"fa",x"f9",x"ff",x"ff",x"fe",x"f9",x"f9",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f5",x"fa",x"f5",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"84",x"88",x"ac",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"d1",x"ad",x"8d",x"8d",x"8d",x"8d",x"ad",x"ad",x"ad",x"ad",x"8d",x"8d",x"8d",x"89",x"89",x"89",x"69",x"8d",x"f5",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"d2",x"ca",x"c6",x"c6",x"ca",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"c6",x"c6",x"ca",x"ca",x"c6",x"ca",x"ee",x"ee",x"c9",x"c6",x"c6",x"c6",x"ca",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ce",x"ca",x"c5",x"c5",x"ca",x"ca",x"ca",x"ca",x"ca",x"c6",x"c5",x"c5",x"ca",x"ca",x"ca",x"c9",x"ca",x"f2",x"c9",x"c9",x"c9",x"c9",x"c9",x"ca",x"ca",x"ca",x"ca",x"ea",x"ea",x"ea",x"ca",x"c6",x"c5",x"c6",x"c9",x"ee",x"ee",x"ca",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"a5",x"c5",x"c6",x"c6",x"c6",x"c9",x"cd",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d5",x"fa",x"fa",x"fa",x"fa",x"fa",x"ff",x"ff",x"fe",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"fe",x"f5",x"f1",x"f5",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f5",x"f1",x"f5",x"d1",x"4d",x"0d",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"31",x"31",x"2d",x"2d",x"2d",x"4d",x"51",x"31",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2c",x"51",x"71",x"b6",x"da",x"da",x"fb",x"fb",x"d6",x"d6",x"b6",x"71",x"2d",x"4d",x"b1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"ac",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"a8",x"f6",x"fa",x"f5",x"fa",x"ff",x"ff",x"fe",x"f5",x"f9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"d1",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"ac",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"d5",x"ad",x"89",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"89",x"89",x"89",x"69",x"89",x"d5",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f2",x"c6",x"a6",x"c6",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"ca",x"f2",x"ca",x"c5",x"c6",x"c6",x"c6",x"ca",x"ea",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"ca",x"c5",x"c5",x"c6",x"c6",x"ca",x"ca",x"c6",x"c6",x"c5",x"c6",x"ca",x"ce",x"ca",x"c6",x"c5",x"ea",x"ee",x"ca",x"c9",x"c9",x"c9",x"ca",x"ca",x"c9",x"c5",x"c5",x"ca",x"ea",x"ea",x"ca",x"c5",x"c5",x"ca",x"ee",x"ee",x"ca",x"a6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"a5",x"c6",x"c6",x"c5",x"cd",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f1",x"d5",x"fb",x"ff",x"fa",x"f5",x"f5",x"fa",x"fa",x"ff",x"ff",x"ff",x"fa",x"fa",x"fe",x"f9",x"f5",x"ff",x"fa",x"f1",x"f1",x"f1",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f1",x"f5",x"f5",x"d1",x"6d",x"2d",x"09",x"09",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"0c",x"71",x"b6",x"da",x"db",x"db",x"da",x"db",x"db",x"d6",x"d6",x"d6",x"b6",x"b2",x"b2",x"d5",x"f5",x"f5",x"f1",x"f1",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"ac",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"b1",x"f5",x"f9",x"fe",x"ff",x"ff",x"fe",x"f5",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"fe",x"fe",x"fe",x"fe",x"f5",x"a8",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"84",x"64",x"88",x"ac",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"d5",x"b1",x"8d",x"89",x"69",x"89",x"89",x"89",x"89",x"69",x"69",x"69",x"89",x"ad",x"d5",x"f9",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f2",x"ce",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"ca",x"ca",x"ee",x"ee",x"ca",x"c5",x"c5",x"c6",x"c6",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c5",x"ca",x"ee",x"ca",x"c6",x"c5",x"c9",x"ee",x"ee",x"ca",x"c5",x"c5",x"c6",x"c6",x"c6",x"c5",x"c5",x"c5",x"c5",x"ca",x"ca",x"c9",x"c9",x"ee",x"ee",x"ee",x"cd",x"cd",x"cd",x"cd",x"f1",x"f1",x"cd",x"c9",x"c6",x"c6",x"a5",x"a5",x"a6",x"c6",x"cd",x"d1",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f5",x"f5",x"fa",x"ff",x"ff",x"fa",x"fa",x"f5",x"f5",x"fa",x"ff",x"ff",x"f5",x"f5",x"fe",x"ff",x"fa",x"f5",x"fa",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5"),
(x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"d1",x"8d",x"4d",x"09",x"09",x"09",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"0d",x"51",x"b6",x"db",x"fb",x"db",x"db",x"db",x"db",x"da",x"d6",x"d6",x"d6",x"d6",x"d6",x"b6",x"d6",x"d5",x"f1",x"f1",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f1",x"f5",x"f5",x"d1",x"ac",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"f5",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fa",x"f9",x"fa",x"fe",x"fe",x"fa",x"ad",x"84",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"ac",x"ac",x"d1",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"d6",x"d1",x"b1",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"ad",x"b1",x"d5",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f6",x"d2",x"ce",x"c9",x"c9",x"c9",x"c9",x"ca",x"c6",x"c6",x"a6",x"c6",x"c6",x"c6",x"c6",x"ca",x"ee",x"ee",x"c9",x"c9",x"ca",x"c6",x"ca",x"ca",x"ca",x"ca",x"ca",x"c6",x"c5",x"c5",x"c5",x"c5",x"c6",x"c6",x"c5",x"c6",x"ca",x"c9",x"ea",x"ea",x"c6",x"c6",x"cd",x"f1",x"ee",x"ee",x"ea",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c9",x"ca",x"ca",x"ca",x"ca",x"c9",x"ee",x"ee",x"ee",x"ce",x"d1",x"d5",x"f1",x"f5",x"f5",x"f5",x"f5",x"d1",x"cd",x"cd",x"cd",x"cd",x"cd",x"cd",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f6",x"fa",x"fe",x"ff",x"fa",x"fa",x"f5",x"f5",x"fa",x"fe",x"fe",x"f5",x"f5",x"fa",x"fe",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f5",x"f5",x"f5",x"d1",x"6d",x"09",x"09",x"09",x"09",x"09",x"0d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"09",x"2d",x"da",x"fb",x"db",x"da",x"db",x"db",x"ff",x"fb",x"da",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"96",x"92",x"d1",x"f5",x"f5",x"f9",x"f9",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"cd",x"88",x"88",x"88",x"88",x"88",x"88",x"f5",x"fe",x"fe",x"fa",x"f9",x"f5",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fa",x"f9",x"f9",x"fe",x"fe",x"fa",x"d1",x"84",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"a8",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"b1",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"fa",x"fa",x"f5",x"d5",x"d5",x"b1",x"d1",x"d5",x"d5",x"f9",x"f9",x"f9",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f5",x"d1",x"cd",x"ce",x"ce",x"ca",x"c5",x"c5",x"a5",x"c6",x"c6",x"c6",x"c6",x"c5",x"ea",x"ee",x"ee",x"ee",x"ea",x"ca",x"ca",x"c6",x"c6",x"c6",x"c6",x"c6",x"c5",x"c5",x"c5",x"c6",x"c5",x"c5",x"c9",x"ca",x"ee",x"ee",x"ca",x"c6",x"cd",x"f5",x"f5",x"ea",x"f2",x"f2",x"ee",x"ee",x"ce",x"ce",x"ee",x"ee",x"cd",x"ee",x"ee",x"ee",x"ee",x"ee",x"ee",x"c6",x"a6",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"fa",x"fb",x"f5",x"fe",x"ff",x"d5",x"f5",x"fa",x"fa",x"f5",x"f5",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"d1",x"b1",x"6d",x"4d",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"0d",x"0d",x"0d",x"0d",x"09",x"09",x"4d",x"b6",x"db",x"da",x"db",x"db",x"db",x"db",x"db",x"db",x"d6",x"d6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"b2",x"b2",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"d1",x"d1",x"ac",x"88",x"84",x"84",x"f5",x"fe",x"fa",x"f9",x"f5",x"f5",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"f9",x"f5",x"f9",x"fa",x"fa",x"f9",x"f5",x"ac",x"88",x"88",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"84",x"84",x"88",x"a8",x"ad",x"d1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"fa",x"f9",x"f9",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"d1",x"d1",x"d2",x"f1",x"f1",x"ca",x"c5",x"ca",x"ea",x"ea",x"ca",x"ca",x"ea",x"ea",x"ee",x"e9",x"e9",x"ca",x"ca",x"c9",x"ea",x"ea",x"ea",x"ea",x"ca",x"ea",x"ea",x"ca",x"c6",x"c6",x"d1",x"f9",x"f5",x"c9",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"ea",x"c6",x"cd",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f5",x"d5",x"fe",x"ff",x"f1",x"fa",x"fe",x"d5",x"f5",x"f9",x"f1",x"ec",x"f4",x"fa",x"f6",x"f5",x"f5",x"f9",x"f5",x"d1",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"d1",x"91",x"6d",x"4d",x"2d",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"08",x"2d",x"96",x"fb",x"db",x"da",x"da",x"da",x"d6",x"d6",x"d6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b2",x"92",x"91",x"92",x"91",x"b1",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"ac",x"a8",x"88",x"f5",x"fa",x"fa",x"f5",x"f5",x"f5",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"f5",x"fa",x"fa",x"f9",x"f5",x"f5",x"d1",x"88",x"88",x"a8",x"a8",x"a8",x"88",x"88",x"88",x"88",x"a8",x"a8",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"a8",x"ac",x"d1",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f1",x"c9",x"c6",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c9",x"c9",x"e9",x"ea",x"ea",x"ca",x"ea",x"ea",x"ea",x"ea",x"ea",x"ca",x"ca",x"c6",x"c6",x"cd",x"f5",x"f9",x"f5",x"ed",x"c6",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"ca",x"c6",x"c6",x"ca",x"ca",x"c6",x"c9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"d5",x"d5",x"fa",x"fe",x"d1",x"f5",x"fa",x"d5",x"f5",x"f9",x"f1",x"ec",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"f1",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"d1",x"f5",x"f5",x"f5",x"f5",x"d1",x"b1",x"6d",x"4d",x"2d",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"29",x"92",x"fb",x"ff",x"db",x"db",x"d6",x"b6",x"d6",x"da",x"d6",x"d6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b2",x"92",x"91",x"91",x"6d",x"72",x"d6",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"f5",x"fa",x"fa",x"f5",x"f5",x"fa",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"ff",x"ff",x"fa",x"ff",x"fe",x"f9",x"f5",x"f5",x"d1",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"84",x"84",x"88",x"ac",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f5",x"f5",x"fa",x"f5",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"d1",x"c9",x"c6",x"c6",x"ca",x"a6",x"a5",x"a5",x"a5",x"a5",x"c6",x"c6",x"c6",x"ca",x"ca",x"ca",x"c6",x"c6",x"c6",x"c6",x"c6",x"c6",x"c9",x"d5",x"f9",x"f5",x"f5",x"f5",x"c5",x"ca",x"ca",x"c5",x"c5",x"c6",x"c6",x"c6",x"c5",x"c5",x"c5",x"c6",x"c6",x"c6",x"a6",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d1",x"d1",x"f9",x"d1",x"f0",x"f5",x"d5",x"d5",x"fa",x"f9",x"f5",x"f5",x"f5",x"fa",x"f5",x"f5",x"d1",x"d1",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f1",x"d1",x"d1",x"b1",x"91",x"91",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"91",x"91",x"ad",x"b1",x"b6",x"db",x"fb",x"fb",x"fb",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b2",x"92",x"92",x"91",x"6d",x"92",x"b2",x"b6",x"b6",x"92",x"91",x"d5",x"f9",x"f5",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"fe",x"fe",x"ff",x"ff",x"ff",x"fe",x"fa",x"fa",x"fe",x"fe",x"ff",x"fe",x"fa",x"f9",x"f5",x"f5",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"84",x"84",x"84",x"88",x"88",x"ac",x"ad",x"d1",x"d1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"f9",x"f5",x"f5",x"f5",x"f9",x"f5",x"f1",x"cd",x"c6",x"a6",x"c6",x"a5",x"c6",x"c6",x"c5",x"c5",x"c6",x"c5",x"c6",x"a6",x"c6",x"a6",x"a6",x"c6",x"a5",x"a6",x"c9",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"c6",x"c6",x"c5",x"c5",x"c6",x"c6",x"c5",x"a5",x"c6",x"c6",x"a6",x"c6",x"c6",x"cd",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"f5",x"f5",x"f0",x"f0",x"f5",x"f5",x"f5",x"d1",x"d1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"d1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"f5",x"f1",x"f5",x"fa",x"db",x"db",x"da",x"db",x"fb",x"ff",x"da",x"da",x"d6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b2",x"b2",x"b2",x"92",x"92",x"b6",x"b6",x"db",x"b6",x"92",x"6d",x"b1",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"fa",x"fe",x"fe",x"ff",x"ff",x"fe",x"fa",x"fa",x"f9",x"f9",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"f5",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"ac",x"ad",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fe",x"fa",x"fa",x"fa",x"fe",x"fe",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"cd",x"c5",x"c6",x"a5",x"c6",x"c6",x"c5",x"a5",x"c6",x"a6",x"c6",x"a5",x"c5",x"c6",x"c5",x"c5",x"c5",x"ca",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"c9",x"c6",x"c6",x"c5",x"c6",x"c6",x"a6",x"c5",x"ce",x"cd",x"c9",x"a6",x"c9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d5",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"cc",x"d0",x"f1",x"d1",x"d1",x"d1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"d1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"d6",x"db",x"db",x"db",x"da",x"da",x"d6",x"db",x"ff",x"ff",x"db",x"d6",x"d6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"91",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d1",x"f5",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"f5",x"f5",x"f5",x"fa",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"ad",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"84",x"84",x"84",x"84",x"88",x"88",x"ac",x"d1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"cd",x"a6",x"a6",x"a6",x"c5",x"a6",x"a6",x"a2",x"ca",x"cd",x"cd",x"cd",x"ce",x"cd",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"cd",x"c6",x"c6",x"c6",x"a6",x"a6",x"cd",x"f5",x"f5",x"d1",x"c9",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"d1",x"d1",x"d1",x"d1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f5",x"d6",x"db",x"db",x"db",x"db",x"db",x"d6",x"da",x"db",x"db",x"da",x"d6",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"8d",x"6d",x"6d",x"6d",x"49",x"6d",x"d5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"d5",x"fa",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"f0",x"f0",x"f9",x"f9",x"f4",x"f0",x"f0",x"f0",x"f5",x"f0",x"ad",x"84",x"84",x"84",x"88",x"88",x"88",x"88",x"a8",x"ac",x"ac",x"ad",x"d1",x"d1",x"d1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f1",x"d1",x"cd",x"cd",x"c9",x"c9",x"cd",x"cd",x"d1",x"d5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"cd",x"cd",x"c9",x"ca",x"cd",x"f5",x"f5",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"d6",x"da",x"db",x"db",x"db",x"db",x"db",x"d6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"91",x"91",x"8d",x"8d",x"8d",x"6d",x"6d",x"6d",x"6d",x"92",x"91",x"d5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f5",x"fe",x"ff",x"fe",x"fa",x"fe",x"fe",x"fe",x"f9",x"f0",x"f4",x"fe",x"f9",x"f5",x"f0",x"ec",x"f0",x"f5",x"f0",x"d1",x"88",x"88",x"88",x"88",x"ac",x"ac",x"ad",x"d1",x"d1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"d1",x"d1",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"d1",x"cd",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"d1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"d6",x"db",x"db",x"db",x"db",x"da",x"d6",x"d6",x"d6",x"b6",x"b6",x"b6",x"92",x"8d",x"92",x"b2",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"91",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"8d",x"d5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f9",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"ff",x"fa",x"f5",x"f0",x"ec",x"f5",x"fa",x"f5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f5",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f5",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"db",x"db",x"db",x"d6",x"b6",x"da",x"d6",x"d6",x"b6",x"b6",x"b6",x"b6",x"b2",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"8d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"49",x"49",x"b1",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"f5",x"fe",x"ff",x"fe",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"f9",x"f5",x"fa",x"fa",x"fa",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"bb",x"db",x"db",x"b6",x"b6",x"d6",x"d6",x"d6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"91",x"6d",x"6d",x"6d",x"91",x"b2",x"91",x"49",x"69",x"25",x"b1",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"d5",x"fa",x"fe",x"fe",x"fe",x"f9",x"f9",x"f9",x"fe",x"ff",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"f9",x"fa",x"d5",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"b6",x"da",x"da",x"d6",x"d6",x"d6",x"d6",x"b6",x"d6",x"b6",x"b6",x"b6",x"b6",x"b2",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"6d",x"6d",x"6d",x"92",x"b2",x"8d",x"69",x"69",x"69",x"25",x"8d",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"d1",x"f5",x"f5",x"d5",x"fa",x"fe",x"fa",x"fe",x"f9",x"f9",x"f5",x"f9",x"fa",x"f5",x"f4",x"f0",x"ec",x"f1",x"f5",x"f5",x"f0",x"f1",x"f5",x"d1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d6",x"b6",x"b6",x"d6",x"da",x"d6",x"d6",x"b6",x"b6",x"b6",x"b6",x"b2",x"b2",x"b2",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"29",x"8d",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"d5",x"fa",x"fa",x"fa",x"fa",x"f5",x"f4",x"f5",x"fa",x"f5",x"f0",x"ec",x"ec",x"f0",x"f5",x"f0",x"f0",x"f1",x"d5",x"d1",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"92",x"b6",x"b6",x"d6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b2",x"b2",x"b2",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"8d",x"6d",x"6d",x"6d",x"92",x"b2",x"91",x"69",x"49",x"69",x"49",x"49",x"29",x"8d",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"d1",x"d1",x"f5",x"f9",x"f9",x"fe",x"f5",x"f0",x"f9",x"fe",x"f5",x"f0",x"ec",x"ec",x"f5",x"f5",x"f0",x"f0",x"f5",x"d1",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"fe",x"fe",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fe",x"fe",x"fe",x"fa",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b2",x"92",x"b2",x"92",x"92",x"91",x"91",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"6d",x"6d",x"69",x"69",x"49",x"49",x"49",x"49",x"b1",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d1",x"d1",x"f9",x"f5",x"f5",x"f9",x"f5",x"fa",x"fa",x"fa",x"fa",x"f9",x"f5",x"fa",x"fa",x"f9",x"fa",x"f6",x"d1",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"ff",x"ff",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"92",x"92",x"92",x"92",x"92",x"b2",x"b2",x"b2",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"8d",x"6d",x"6d",x"8d",x"91",x"92",x"92",x"92",x"6d",x"69",x"69",x"69",x"49",x"49",x"49",x"49",x"6d",x"d1",x"f5",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d1",x"d1",x"f5",x"f4",x"f4",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"fa",x"fa",x"f9",x"f9",x"f9",x"d5",x"d1",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"91",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b2",x"92",x"8d",x"69",x"69",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"d1",x"f5",x"f5",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"d1",x"ad",x"f0",x"f0",x"f5",x"f5",x"f4",x"f0",x"f0",x"ec",x"f0",x"fa",x"f9",x"f5",x"f5",x"f5",x"d1",x"d5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fe",x"fe",x"fe",x"ff",x"ff",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"f9",x"f9",x"f9",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"d1",x"92",x"92",x"b2",x"b6",x"96",x"92",x"92",x"92",x"92",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"49",x"49",x"29",x"69",x"b1",x"f1",x"f5",x"f5",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f1",x"d1",x"d1",x"d0",x"f5",x"f5",x"f0",x"f0",x"f0",x"ec",x"f0",x"f9",x"f5",x"d0",x"d1",x"d1",x"d1",x"f1",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fa",x"da",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"b1",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"6d",x"6d",x"49",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"b1",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f1",x"d1",x"d1",x"d5",x"f5",x"f0",x"f0",x"f0",x"ec",x"d0",x"f5",x"d1",x"d1",x"d1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fa",x"da",x"da",x"da",x"d5",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"d1",x"91",x"6d",x"6d",x"8d",x"92",x"92",x"b2",x"92",x"92",x"92",x"92",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"8d",x"d1",x"f5",x"f1",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f1",x"f5",x"f1",x"d1",x"d1",x"b1",x"d1",x"d1",x"d1",x"d1",x"b1",x"d1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fe",x"ff",x"ff",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"d5",x"d1",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"d1",x"b1",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"8d",x"b1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f5",x"da",x"ff",x"ff",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"d6",x"b1",x"d5",x"f5",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d1",x"b1",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"8d",x"d1",x"f5",x"f5",x"f5",x"f1",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"f9",x"f5",x"d5",x"fa",x"fa",x"fa",x"fa",x"da",x"da",x"da",x"d5",x"d1",x"b1",x"d5",x"f5",x"f9",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"f9",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f1",x"f5",x"f5",x"f5",x"b1",x"8d",x"6d",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"8d",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"f9",x"f5",x"d5",x"b1",x"d6",x"d6",x"d5",x"b5",x"b1",x"b1",x"b1",x"d1",x"d5",x"f5",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"f9",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d1",x"d1",x"b1",x"91",x"8d",x"8d",x"6d",x"6d",x"6d",x"8d",x"8d",x"b1",x"b1",x"d1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f5",x"d1",x"d1",x"d1",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"f5",x"f5",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"da",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d1",x"b1",x"b1",x"b1",x"b1",x"d1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f5",x"d1",x"d1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"d6",x"d6",x"d6",x"d6",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"ff",x"fe",x"d6",x"d6",x"d6",x"d5",x"d6",x"d5",x"da",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fa",x"da",x"da",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"ff",x"ff",x"ff",x"fe",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d6",x"d5",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"d6",x"fa",x"fe",x"ff",x"ff",x"ff",x"fe",x"ff",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d6",x"d1",x"d1",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"fe",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f5",x"d6",x"da",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fa",x"fa",x"da",x"d6",x"d6",x"fa",x"fa",x"fa",x"d6",x"d5",x"d5",x"d1",x"b1",x"d1",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"d5",x"d6",x"d6",x"fa",x"fa",x"fa",x"fa",x"fa",x"da",x"d6",x"d6",x"d5",x"d5",x"d5",x"d6",x"d6",x"d5",x"d5",x"d5",x"b1",x"b1",x"b1",x"d5",x"f9",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"d5",x"d6",x"d6",x"d5",x"d6",x"d6",x"d6",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d1",x"d1",x"b1",x"b1",x"d1",x"f5",x"f5",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f5",x"d5",x"d5",x"d6",x"d6",x"d6",x"d6",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"b1",x"b1",x"b1",x"d1",x"d5",x"f5",x"f5",x"f5",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f5",x"d5",x"d1",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d1",x"b1",x"b1",x"b1",x"d1",x"d1",x"d1",x"d1",x"f5",x"f5",x"f5",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"fa",x"f9",x"f5",x"f5",x"d5",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"fa",x"f9",x"f9",x"f5",x"d5",x"d5",x"d5",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d1",x"d5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d1",x"d1",x"d1",x"d1",x"d1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"fa",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5"),
(x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1"),
(x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1"),
(x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1"),
(x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1"),
(x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1"),
(x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1"),
(x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1"),
(x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f5",x"f1",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1"),
(x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1"),
(x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1")
);

begin

process ( RESETn, CLK)
begin
    if RESETn = '0' then
        mVGA_RGB	<=  (others => '0') ; 	
    	drawing_request	<=  '0' ;
	elsif rising_edge(CLK) then
		mVGA_RGB	<=  object_color(oCoord_X, oCoord_Y);
		drawing_request	<= '1';
	end if;

end process;

		
end behav;		
