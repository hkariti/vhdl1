--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity QubeTable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end QubeTable;

architecture arch of QubeTable is
constant array_size 			: integer := 256 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal Qube_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant Qube_table : table_type := (
---start 0 v
X"C180",
X"C2F5",
X"C463",
X"C5CB",
X"C72E",
X"C88B",
X"C9E3",
X"CB35",
X"CC81",
X"CDC8",
X"CF09",
X"D045",
X"D17C",
X"D2AD",
X"D3D9",
X"D500",
X"D622",
X"D73E",
X"D856",
X"D968",
X"DA76",
X"DB7E",
X"DC82",
X"DD81",
X"DE7A",
X"DF70",
X"E060",
X"E14C",
X"E233",
X"E316",
X"E3F4",
X"E4CD",
X"E5A2",
X"E673",
X"E740",
X"E808",
X"E8CC",
X"E98B",
X"EA47",
X"EAFE",
X"EBB1",
X"EC61",
X"ED0C",
X"EDB3",
X"EE57",
X"EEF6",
X"EF92",
X"F02A",
X"F0BE",
X"F14F",
X"F1DC",
X"F265",
X"F2EB",
X"F36E",
X"F3ED",
X"F469",
X"F4E1",
X"F556",
X"F5C8",
X"F636",
X"F6A2",
X"F70A",
X"F76F",
X"F7D1",
X"F830",
X"F88D",
X"F8E6",
X"F93D",
X"F991",
X"F9E2",
X"FA30",
X"FA7C",
X"FAC5",
X"FB0B",
X"FB4F",
X"FB91",
X"FBD0",
X"FC0C",
X"FC47",
X"FC7F",
X"FCB5",
X"FCE8",
X"FD1A",
X"FD49",
X"FD77",
X"FDA2",
X"FDCB",
X"FDF3",
X"FE18",
X"FE3C",
X"FE5E",
X"FE7E",
X"FE9D",
X"FEB9",
X"FED5",
X"FEEE",
X"FF06",
X"FF1D",
X"FF33",
X"FF46",
X"FF59",
X"FF6A",
X"FF7A",
X"FF89",
X"FF97",
X"FFA4",
X"FFAF",
X"FFBA",
X"FFC3",
X"FFCC",
X"FFD4",
X"FFDB",
X"FFE1",
X"FFE7",
X"FFEC",
X"FFF0",
X"FFF3",
X"FFF6",
X"FFF9",
X"FFFB",
X"FFFD",
X"FFFE",
X"FFFF",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0001",
X"0002",
X"0003",
X"0005",
X"0007",
X"000A",
X"000D",
X"0010",
X"0014",
X"0019",
X"001F",
X"0025",
X"002C",
X"0034",
X"003D",
X"0046",
X"0051",
X"005C",
X"0069",
X"0077",
X"0086",
X"0096",
X"00A7",
X"00BA",
X"00CD",
X"00E3",
X"00FA",
X"0112",
X"012B",
X"0147",
X"0163",
X"0182",
X"01A2",
X"01C4",
X"01E8",
X"020D",
X"0235",
X"025E",
X"0289",
X"02B7",
X"02E6",
X"0318",
X"034B",
X"0381",
X"03B9",
X"03F4",
X"0430",
X"046F",
X"04B1",
X"04F5",
X"053B",
X"0584",
X"05D0",
X"061E",
X"066F",
X"06C3",
X"071A",
X"0773",
X"07D0",
X"082F",
X"0891",
X"08F6",
X"095E",
X"09CA",
X"0A38",
X"0AAA",
X"0B1F",
X"0B97",
X"0C13",
X"0C92",
X"0D15",
X"0D9B",
X"0E24",
X"0EB1",
X"0F42",
X"0FD6",
X"106E",
X"110A",
X"11A9",
X"124D",
X"12F4",
X"139F",
X"144F",
X"1502",
X"15B9",
X"1675",
X"1734",
X"17F8",
X"18C0",
X"198D",
X"1A5E",
X"1B33",
X"1C0C",
X"1CEA",
X"1DCD",
X"1EB4",
X"1FA0",
X"2090",
X"2186",
X"227F",
X"237E",
X"2482",
X"258A",
X"2698",
X"27AA",
X"28C2",
X"29DE",
X"2B00",
X"2C27",
X"2D53",
X"2E84",
X"2FBB",
X"30F7",
X"3238",
X"337F",
X"34CB",
X"361D",
X"3775",
X"38D2",
X"3A35",
X"3B9D",
X"3D0B"
 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= Qube_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;